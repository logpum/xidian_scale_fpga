
//
// Verific Verilog Description of module T35_Sensor_DDR3_LCD_Test
//

module T35_Sensor_DDR3_LCD_Test (Axi_Clk, tx_slowclk, tx_fastclk, pll_clk_200m, 
            hdmi_clk1x_i, hdmi_clk2x_i, hdmi_clk5x_i, PllLocked, DdrCtrl_CFG_RST_N, 
            DdrCtrl_CFG_SEQ_RST, DdrCtrl_CFG_SEQ_START, DdrCtrl_AID_0, 
            DdrCtrl_AADDR_0, DdrCtrl_ALEN_0, DdrCtrl_ASIZE_0, DdrCtrl_ABURST_0, 
            DdrCtrl_ALOCK_0, DdrCtrl_AVALID_0, DdrCtrl_AREADY_0, DdrCtrl_ATYPE_0, 
            DdrCtrl_WID_0, DdrCtrl_WDATA_0, DdrCtrl_WSTRB_0, DdrCtrl_WLAST_0, 
            DdrCtrl_WVALID_0, DdrCtrl_WREADY_0, DdrCtrl_RID_0, DdrCtrl_RDATA_0, 
            DdrCtrl_RLAST_0, DdrCtrl_RVALID_0, DdrCtrl_RREADY_0, DdrCtrl_RRESP_0, 
            DdrCtrl_BID_0, DdrCtrl_BVALID_0, DdrCtrl_BREADY_0, LED, 
            cmos_sclk, cmos_sdat_IN, cmos_sdat_OUT, cmos_sdat_OE, cmos_pclk, 
            cmos_vsync, cmos_href, cmos_data, cmos_ctl0, cmos_ctl1, 
            cmos_ctl2, cmos_ctl3, hdmi_tx0_o, hdmi_tx1_o, hdmi_tx2_o, 
            hdmi_txc_o, lcd_pwm, lvds_tx_clk_DATA, lvds_tx0_DATA, lvds_tx1_DATA, 
            lvds_tx2_DATA, lvds_tx3_DATA, jtag_inst1_CAPTURE, jtag_inst1_DRCK, 
            jtag_inst1_RESET, jtag_inst1_RUNTEST, jtag_inst1_SEL, jtag_inst1_SHIFT, 
            jtag_inst1_TCK, jtag_inst1_TDI, jtag_inst1_TMS, jtag_inst1_UPDATE, 
            jtag_inst1_TDO);
    input Axi_Clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input tx_slowclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input tx_fastclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input pll_clk_200m /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input hdmi_clk1x_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input hdmi_clk2x_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input hdmi_clk5x_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [1:0]PllLocked /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_CFG_RST_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_CFG_SEQ_RST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_CFG_SEQ_START /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_AID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [31:0]DdrCtrl_AADDR_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_ALEN_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [2:0]DdrCtrl_ASIZE_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]DdrCtrl_ABURST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]DdrCtrl_ALOCK_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_AVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input DdrCtrl_AREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_ATYPE_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_WID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [127:0]DdrCtrl_WDATA_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [15:0]DdrCtrl_WSTRB_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_WLAST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_WVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input DdrCtrl_WREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]DdrCtrl_RID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [127:0]DdrCtrl_RDATA_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_RLAST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_RVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_RREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [1:0]DdrCtrl_RRESP_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]DdrCtrl_BID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_BVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_BREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]LED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output cmos_sclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input cmos_sdat_IN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output cmos_sdat_OUT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output cmos_sdat_OE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input cmos_pclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input cmos_vsync /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input cmos_href /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]cmos_data /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output cmos_ctl0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input cmos_ctl1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output cmos_ctl2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output cmos_ctl3 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_tx0_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_tx1_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_tx2_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_txc_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output lcd_pwm /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx_clk_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx0_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx1_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx2_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx3_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input jtag_inst1_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst1_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    wire \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire n592_2;
    wire n603_2;
    wire n614_2;
    wire n9_2;
    wire \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire n602_2;
    wire n601_2;
    wire n600_2;
    wire n599_2;
    
    wire n186, n187, \ResetShiftReg[0] , \Axi0ResetReg[0] , r_hdmi_rst_n, 
        rc_hdmi_tx, \PowerOnResetCnt[0] , \ResetShiftReg[1] , \Axi0ResetReg[1] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] , \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] , n205, n206, \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] , n228, n229, \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] , 
        n231, n232, \u_i2c_timing_ctrl_16reg_16bit/current_state[0] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk , \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en , 
        \i2c_config_index[0] , \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0] , \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5 , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4 , \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3 , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2 , \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1 , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_ack , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15] , 
        \u_i2c_timing_ctrl_16reg_16bit/current_state[1] , \u_i2c_timing_ctrl_16reg_16bit/current_state[2] , 
        \u_i2c_timing_ctrl_16reg_16bit/current_state[3] , \u_i2c_timing_ctrl_16reg_16bit/current_state[4] , 
        \i2c_config_index[1] , \i2c_config_index[2] , \i2c_config_index[3] , 
        \i2c_config_index[4] , \i2c_config_index[5] , \i2c_config_index[6] , 
        \i2c_config_index[7] , \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] , \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] , \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3] , \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5] , \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19] , n345, n346, n347, 
        n348, n349, n350, n351, n352, n353, n354, n355, n356, 
        n357, n358, n359, n360, n361, n362, n363, n364, n365, 
        n366, n367, n368, n369, n370, n371, n372, n373, n374, 
        n375, n376, n377, n378, n379, n380, n381, n382, n383, 
        n384, n385, n386, n387, n388, n389, n390, n391, n392, 
        n393, n394, n395, n396, n397, n398, n399, n400, n401, 
        n402, n403, n404, n405, n406, n407, n408, n409, n410, 
        n411, n412, n413, n414, n415, n416, n417, n418, n419, 
        n420, n421, n422, n423, n424, n425, n426, n427, n428, 
        n429, n430, n431, n432, n433, n434, n435, n436, n437, 
        n438, n439, n440, \u_CMOS_Capture_RAW_Gray/cmos_href_r[0] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0] , \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0] , 
        n445, n446, \u_CMOS_Capture_RAW_Gray/line_cnt[0] , \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] , 
        \u_CMOS_Capture_RAW_Gray/frame_sync_flag , n453, n454, n455, 
        n461, n462, \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] , \u_CMOS_Capture_RAW_Gray/cmos_href_r[1] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1] , \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3] , \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5] , \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7] , \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2] , \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4] , \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6] , \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[1] , \u_CMOS_Capture_RAW_Gray/line_cnt[2] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[3] , \u_CMOS_Capture_RAW_Gray/line_cnt[4] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[5] , \u_CMOS_Capture_RAW_Gray/line_cnt[6] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[7] , \u_CMOS_Capture_RAW_Gray/line_cnt[8] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[9] , \u_CMOS_Capture_RAW_Gray/line_cnt[10] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[11] , \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] , 
        n531, n532, n541, n542, n543, n544, n545, n546, n547, 
        n548, n549, n550, n551, n552, n553, n554, n555, n556, 
        n557, n558, n559, n560, n561, n562, n563, n564, n565, 
        n566, n567, n568, \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1] , 
        n575, n576, n600, n601, n602, \u_sensor_frame_count/cmos_fps_cnt[0] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n105 , \u_sensor_frame_count/cmos_vsync_r[0] , 
        \u_sensor_frame_count/delay_cnt[0] , \u_sensor_frame_count/delay_cnt[1] , 
        \u_sensor_frame_count/delay_cnt[2] , \u_sensor_frame_count/delay_cnt[3] , 
        \u_sensor_frame_count/delay_cnt[4] , \u_sensor_frame_count/delay_cnt[5] , 
        \u_sensor_frame_count/delay_cnt[6] , \u_sensor_frame_count/delay_cnt[7] , 
        \u_sensor_frame_count/delay_cnt[8] , \u_sensor_frame_count/delay_cnt[9] , 
        \u_sensor_frame_count/delay_cnt[10] , \u_sensor_frame_count/delay_cnt[11] , 
        \u_sensor_frame_count/delay_cnt[12] , \u_sensor_frame_count/delay_cnt[13] , 
        \u_sensor_frame_count/delay_cnt[14] , \u_sensor_frame_count/delay_cnt[15] , 
        \u_sensor_frame_count/delay_cnt[16] , \u_sensor_frame_count/delay_cnt[17] , 
        \u_sensor_frame_count/delay_cnt[18] , \u_sensor_frame_count/delay_cnt[19] , 
        \u_sensor_frame_count/delay_cnt[20] , \u_sensor_frame_count/delay_cnt[21] , 
        \u_sensor_frame_count/delay_cnt[22] , \u_sensor_frame_count/delay_cnt[23] , 
        \u_sensor_frame_count/delay_cnt[24] , \u_sensor_frame_count/delay_cnt[25] , 
        \u_sensor_frame_count/delay_cnt[26] , \u_sensor_frame_count/delay_cnt[27] , 
        n636, \u_sensor_frame_count/cmos_fps_cnt[2] , \u_sensor_frame_count/cmos_fps_cnt[3] , 
        \u_sensor_frame_count/cmos_fps_cnt[4] , \u_sensor_frame_count/cmos_fps_cnt[5] , 
        \u_sensor_frame_count/cmos_fps_cnt[6] , \u_sensor_frame_count/cmos_fps_cnt[7] , 
        \u_sensor_frame_count/cmos_fps_cnt[8] , n646, n648, n650, n651, 
        n652, n653, n654, n655, n656, n657, n658, n659, n660, 
        n661, n662, n663, n664, n665, n666, n667, n668, n669, 
        n670, n671, n672, n673, n674, n675, n676, n677, n678, 
        n679, n680, \u_sensor_frame_count/cmos_vsync_r[1] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 , 
        n693, n694, n695, n696, n697, \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n98 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n99 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n102 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n104 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n96 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n93 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n90 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n87 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n84 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n101 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n95 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n92 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n89 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n86 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n83 , 
        n713, n714, \u_afifo_buf/u_efx_fifo_top/waddr[0] , empty, n717, 
        n718, n719, n720, \u_afifo_buf/u_efx_fifo_top/raddr[0] , n722, 
        n723, n724, n725, n726, n727, \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[1] , \u_afifo_buf/u_efx_fifo_top/waddr[2] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[3] , \u_afifo_buf/u_efx_fifo_top/waddr[4] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[5] , \u_afifo_buf/u_efx_fifo_top/waddr[6] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[7] , \u_afifo_buf/u_efx_fifo_top/waddr[8] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[9] , \u_afifo_buf/u_efx_fifo_top/waddr[10] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[11] , \u_afifo_buf/u_efx_fifo_top/waddr[12] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] , n745, 
        n746, n747, n748, n749, n750, n751, n752, n753, n754, 
        n755, n756, \u_afifo_buf/u_efx_fifo_top/raddr[1] , \u_afifo_buf/u_efx_fifo_top/raddr[2] , 
        \u_afifo_buf/u_efx_fifo_top/raddr[3] , \u_afifo_buf/u_efx_fifo_top/raddr[4] , 
        \u_afifo_buf/u_efx_fifo_top/raddr[5] , \u_afifo_buf/u_efx_fifo_top/raddr[6] , 
        \u_afifo_buf/u_efx_fifo_top/raddr[7] , \u_afifo_buf/u_efx_fifo_top/raddr[8] , 
        \u_afifo_buf/u_efx_fifo_top/raddr[9] , \u_afifo_buf/u_efx_fifo_top/raddr[10] , 
        \u_afifo_buf/u_efx_fifo_top/raddr[11] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] , 
        n777, n778, n779, n780, n781, n782, n783, n784, n785, 
        n786, n787, n788, n789, n790, n791, n792, n793, n794, 
        n795, n796, n797, n798, n799, n800, n801, n802, n803, 
        n804, n805, n806, n807, n808, n809, n810, n811, n812, 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13] , 
        \u_scaler_gray/vs_cnt[0] , n910, n911, tvsync_o, \u_scaler_gray/tvalid_o_r , 
        n914, n915, n916, n917, n918, n919, \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] , 
        n921, n922, n923, n924, n925, n926, \u_scaler_gray/u0_data_stream_ctr/w_addra[0] , 
        n928, n929, n930, n931, \u_scaler_gray/u0_data_stream_ctr/scaler_st[0] , 
        n933, n934, n935, n936, n937, n938, n939, \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0] , 
        \u_scaler_gray/destx[0] , n942, n943, n944, n945, n946, 
        n947, n948, n949, \u_scaler_gray/desty[0] , n951, n952, 
        n954, n955, n956, n957, n958, n959, n960, n961, n962, 
        n963, \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0] , 
        n966, n967, \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0] , 
        \u_scaler_gray/tdata00[0] , \u_scaler_gray/tdata01[0] , \u_scaler_gray/tdata10[0] , 
        \u_scaler_gray/tdata11[0] , n973, n974, n975, n976, \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] , n1010, n1011, 
        n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
        n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
        n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, 
        n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
        n1044, n1045, n1046, n1047, \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[12] , \u_scaler_gray/u0_data_stream_ctr/w_addra[13] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[14] , \u_scaler_gray/u0_data_stream_ctr/w_addra[15] , 
        n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
        n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, 
        n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
        n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
        n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
        n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, 
        \u_scaler_gray/u0_data_stream_ctr/scaler_st[1] , \u_scaler_gray/u0_data_stream_ctr/scaler_st[2] , 
        n1113, n1114, n1115, n1116, \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1] , 
        \u_scaler_gray/destx[1] , \u_scaler_gray/destx[2] , \u_scaler_gray/destx[3] , 
        \u_scaler_gray/destx[4] , \u_scaler_gray/destx[5] , \u_scaler_gray/destx[6] , 
        \u_scaler_gray/destx[7] , \u_scaler_gray/destx[8] , \u_scaler_gray/destx[9] , 
        \u_scaler_gray/destx[10] , \u_scaler_gray/destx[11] , \u_scaler_gray/destx[12] , 
        \u_scaler_gray/destx[13] , \u_scaler_gray/destx[14] , \u_scaler_gray/destx[15] , 
        n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, 
        n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, 
        n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
        n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
        n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
        n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, 
        n1181, n1182, n1183, \u_scaler_gray/desty[1] , \u_scaler_gray/desty[2] , 
        \u_scaler_gray/desty[3] , \u_scaler_gray/desty[4] , \u_scaler_gray/desty[5] , 
        \u_scaler_gray/desty[6] , \u_scaler_gray/desty[7] , \u_scaler_gray/desty[8] , 
        \u_scaler_gray/desty[9] , \u_scaler_gray/desty[10] , \u_scaler_gray/desty[11] , 
        \u_scaler_gray/desty[12] , \u_scaler_gray/desty[13] , \u_scaler_gray/desty[14] , 
        \u_scaler_gray/desty[15] , n1199, n1200, n1201, n1202, n1203, 
        n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, 
        n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
        n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
        n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
        n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, 
        n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, 
        n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
        n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8] , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10] , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11] , 
        n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
        n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, 
        n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, 
        n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, 
        n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, 
        n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
        n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
        n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
        n1336, n1337, n1338, n1339, n1340, \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2] , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4] , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6] , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8] , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10] , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11] , n1363, n1364, 
        n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8] , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10] , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11] , 
        \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1] , \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2] , 
        \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] , \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4] , 
        \u_scaler_gray/tvalid , \u_scaler_gray/tdata00[1] , \u_scaler_gray/tdata00[2] , 
        \u_scaler_gray/tdata00[3] , \u_scaler_gray/tdata00[4] , \u_scaler_gray/tdata00[5] , 
        \u_scaler_gray/tdata00[6] , \u_scaler_gray/tdata00[7] , \u_scaler_gray/tdata01[1] , 
        \u_scaler_gray/tdata01[2] , \u_scaler_gray/tdata01[3] , \u_scaler_gray/tdata01[4] , 
        \u_scaler_gray/tdata01[5] , \u_scaler_gray/tdata01[6] , \u_scaler_gray/tdata01[7] , 
        \u_scaler_gray/tdata10[1] , \u_scaler_gray/tdata10[2] , \u_scaler_gray/tdata10[3] , 
        \u_scaler_gray/tdata10[4] , \u_scaler_gray/tdata10[5] , \u_scaler_gray/tdata10[6] , 
        \u_scaler_gray/tdata10[7] , \u_scaler_gray/tdata11[1] , \u_scaler_gray/tdata11[2] , 
        \u_scaler_gray/tdata11[3] , \u_scaler_gray/tdata11[4] , \u_scaler_gray/tdata11[5] , 
        \u_scaler_gray/tdata11[6] , \u_scaler_gray/tdata11[7] , n1410, 
        n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, 
        n1419, n1420, \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15] , 
        n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, 
        n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
        n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, 
        n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, 
        n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
        n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, 
        n1511, n1512, n1513, n1514, n1515, n1516, n1517, \u_scaler_gray/vs_cnt[1] , 
        \u_scaler_gray/vs_cnt[2] , \u_scaler_gray/vs_cnt[3] , \u_scaler_gray/vs_cnt[4] , 
        \u_scaler_gray/vs_cnt[5] , \u_scaler_gray/vs_cnt[6] , \u_scaler_gray/vs_cnt[7] , 
        \u_scaler_gray/vs_cnt[8] , \u_scaler_gray/vs_cnt[9] , \u_scaler_gray/vs_cnt[10] , 
        \u_scaler_gray/vs_cnt[11] , \u_scaler_gray/vs_cnt[12] , \u_scaler_gray/vs_cnt[13] , 
        \u_scaler_gray/vs_cnt[14] , \u_scaler_gray/vs_cnt[15] , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[0] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0] , 
        n1535, n1536, n1537, n1538, \u_scaler_gray/u1_bilinear_gray/srcy_fix[0] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[1] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[2] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[3] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[4] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[5] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[6] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[7] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[8] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[9] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[10] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[11] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[12] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[13] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[14] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[15] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[16] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[17] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[18] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[19] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[20] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[21] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[22] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[23] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[24] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[25] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[26] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[27] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27] , 
        \u_scaler_gray/u1_bilinear_gray/srcx_fix[9] , \u_scaler_gray/u1_bilinear_gray/srcx_fix[10] , 
        \u_scaler_gray/u1_bilinear_gray/srcx_fix[11] , \u_scaler_gray/srcx_int[0] , 
        \u_scaler_gray/srcx_int[1] , \u_scaler_gray/srcx_int[2] , \u_scaler_gray/srcx_int[3] , 
        \u_scaler_gray/srcx_int[4] , \u_scaler_gray/srcx_int[5] , \u_scaler_gray/srcx_int[6] , 
        \u_scaler_gray/srcx_int[7] , \u_scaler_gray/srcx_int[8] , \u_scaler_gray/srcx_int[9] , 
        \u_scaler_gray/srcx_int[10] , \u_scaler_gray/srcx_int[11] , \u_scaler_gray/srcx_int[12] , 
        \u_scaler_gray/srcx_int[13] , \u_scaler_gray/srcx_int[14] , \u_scaler_gray/srcx_int[15] , 
        n1654, n1655, n1656, n1657, \u_scaler_gray/u1_bilinear_gray/srcy_fix[1] , 
        \u_scaler_gray/u1_bilinear_gray/srcy_fix[2] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[3] , 
        \u_scaler_gray/u1_bilinear_gray/srcy_fix[4] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[5] , 
        \u_scaler_gray/u1_bilinear_gray/srcy_fix[6] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[7] , 
        \u_scaler_gray/u1_bilinear_gray/srcy_fix[8] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[9] , 
        \u_scaler_gray/u1_bilinear_gray/srcy_fix[10] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[11] , 
        \u_scaler_gray/srcy_int[0] , \u_scaler_gray/srcy_int[1] , \u_scaler_gray/srcy_int[2] , 
        \u_scaler_gray/srcy_int[3] , \u_scaler_gray/srcy_int[4] , \u_scaler_gray/srcy_int[5] , 
        \u_scaler_gray/srcy_int[6] , \u_scaler_gray/srcy_int[7] , \u_scaler_gray/srcy_int[8] , 
        \u_scaler_gray/srcy_int[9] , \u_scaler_gray/srcy_int[10] , \u_scaler_gray/srcy_int[11] , 
        \u_scaler_gray/srcy_int[12] , \u_scaler_gray/srcy_int[13] , \u_scaler_gray/srcy_int[14] , 
        \u_scaler_gray/srcy_int[15] , n1685, n1686, n1687, n1688, 
        n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
        n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, 
        n1705, n1706, n1707, \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0] , 
        n1731, n1732, n1733, n1734, n1735, n1736, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
        n1740, n1741, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11] , 
        n1753, n1754, n1783, n1784, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[11] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[12] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[13] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[14] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[15] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[16] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[17] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[18] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[19] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[20] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[21] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[22] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[23] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[11] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[12] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[13] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[14] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[15] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[16] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[17] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[18] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[19] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[20] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[21] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[22] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[23] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[11] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[12] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[13] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[14] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[15] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[16] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[17] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[18] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[19] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[20] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[21] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[22] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[23] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[11] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[12] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[13] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[14] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[15] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[16] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[17] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[18] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[19] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[20] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[21] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[22] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[23] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0] , 
        n1918, n1919, n1920, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0] , 
        n1922, n1923, n1924, n1925, \tdata_o[0] , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9] , 
        \tdata_o[1] , \tdata_o[2] , \tdata_o[3] , \tdata_o[4] , \tdata_o[5] , 
        \tdata_o[6] , \tdata_o[7] , n2054, n2055, n2056, n2057, 
        n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, 
        n2066, n2067, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[19] , 
        n2091, n2092, n2093, n2094, \u_axi4_ctrl/wframe_vsync_dly[0] , 
        n2096, n2097, n2098, n2099, \u_axi4_ctrl/rframe_vsync_dly[0] , 
        n2102, n2103, \u_axi4_ctrl/wframe_index[0] , n2105, n2106, 
        n2107, n2108, \u_axi4_ctrl/rframe_index[0] , n2110, \u_axi4_ctrl/state[0] , 
        n2112, n2113, n2115, n2116, n2117, n2118, n2119, n2120, 
        n2121, n2122, n2123, n2124, n2125, n2126, n2129, n2130, 
        \u_axi4_ctrl/wdata_cnt_dly[0] , \u_axi4_ctrl/rdata_cnt_dly[1] , 
        \u_axi4_ctrl/rdata_cnt_dly[0] , n2134, n2135, n2136, n2137, 
        n2138, n2139, n2140, n2141, n2142, n2143, \u_axi4_ctrl/rfifo_wenb , 
        \u_axi4_ctrl/rfifo_wdata[0] , n2146, n2147, n2148, n2149, 
        n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
        n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, 
        n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, 
        n2174, n2175, n2176, n2177, n2178, n2179, n2180, \u_axi4_ctrl/wframe_vsync_dly[1] , 
        \u_axi4_ctrl/wframe_vsync_dly[2] , \u_axi4_ctrl/wframe_vsync_dly[3] , 
        n2184, n2185, n2186, n2187, n2188, n2189, n2190, \u_axi4_ctrl/rframe_vsync_dly[1] , 
        \u_axi4_ctrl/rframe_vsync_dly[2] , \u_axi4_ctrl/rframe_vsync_dly[3] , 
        n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, 
        \u_axi4_ctrl/wframe_index[1] , n2322, n2323, n2340, n2341, 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] , \u_axi4_ctrl/wfifo_empty , 
        n2346, n2347, n2348, n2349, n2350, n2351, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] , 
        n2353, n2354, n2355, n2356, n2357, n2358, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] , 
        n2374, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
        n2383, n2384, n2385, n2386, n2387, n2388, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] , 
        n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, 
        n2405, n2406, n2407, n2408, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] , 
        n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, 
        n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, 
        n2504, n2505, n2506, n2516, n2517, n2519, n2520, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] , 
        \u_axi4_ctrl/rfifo_empty , n2523, n2524, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] , 
        n2526, n2527, n2528, n2529, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] , 
        n2533, n2534, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] , 
        n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
        n2551, n2552, n2553, n2554, n2555, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] , 
        n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, 
        n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, 
        n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, 
        n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
        n2600, n2601, n2602, n2603, n2604, n2605, n2606, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] , 
        n2687, n2688, n2689, n2690, n2691, n2692, \u_axi4_ctrl/rframe_index[1] , 
        n2694, n2695, n2696, n2697, \u_axi4_ctrl/state[1] , \u_axi4_ctrl/state[2] , 
        n2700, n2701, n2702, n2703, \u_axi4_ctrl/awaddr[10] , \u_axi4_ctrl/awaddr[11] , 
        \u_axi4_ctrl/awaddr[12] , \u_axi4_ctrl/awaddr[13] , \u_axi4_ctrl/awaddr[14] , 
        \u_axi4_ctrl/awaddr[15] , \u_axi4_ctrl/awaddr[16] , \u_axi4_ctrl/awaddr[17] , 
        \u_axi4_ctrl/awaddr[18] , \u_axi4_ctrl/awaddr[19] , \u_axi4_ctrl/awaddr[20] , 
        \u_axi4_ctrl/awaddr[21] , \u_axi4_ctrl/awaddr[22] , \u_axi4_ctrl/awaddr[23] , 
        n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, 
        n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, 
        n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, 
        n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, 
        n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, 
        n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, 
        n2786, n2787, \u_axi4_ctrl/araddr[10] , \u_axi4_ctrl/araddr[11] , 
        \u_axi4_ctrl/araddr[12] , \u_axi4_ctrl/araddr[13] , \u_axi4_ctrl/araddr[14] , 
        \u_axi4_ctrl/araddr[15] , \u_axi4_ctrl/araddr[16] , \u_axi4_ctrl/araddr[17] , 
        \u_axi4_ctrl/araddr[18] , \u_axi4_ctrl/araddr[19] , \u_axi4_ctrl/araddr[20] , 
        \u_axi4_ctrl/araddr[21] , \u_axi4_ctrl/araddr[22] , \u_axi4_ctrl/araddr[23] , 
        n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, 
        n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, 
        n2818, n2819, n2820, n2821, n2822, n2865, n2866, n2867, 
        n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, 
        n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
        n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, 
        n2892, \u_axi4_ctrl/wdata_cnt_dly[1] , \u_axi4_ctrl/wdata_cnt_dly[2] , 
        \u_axi4_ctrl/wdata_cnt_dly[3] , \u_axi4_ctrl/wdata_cnt_dly[4] , 
        \u_axi4_ctrl/wdata_cnt_dly[5] , \u_axi4_ctrl/wdata_cnt_dly[6] , 
        \u_axi4_ctrl/wdata_cnt_dly[7] , \u_axi4_ctrl/wdata_cnt_dly[8] , 
        \u_axi4_ctrl/rdata_cnt_dly[2] , \u_axi4_ctrl/rdata_cnt_dly[3] , 
        \u_axi4_ctrl/rdata_cnt_dly[4] , \u_axi4_ctrl/rdata_cnt_dly[5] , 
        \u_axi4_ctrl/rdata_cnt_dly[6] , \u_axi4_ctrl/rdata_cnt_dly[7] , 
        \u_axi4_ctrl/rdata_cnt_dly[8] , n2908, n2909, n2910, n2911, 
        \u_axi4_ctrl/rfifo_wdata[1] , \u_axi4_ctrl/rfifo_wdata[2] , \u_axi4_ctrl/rfifo_wdata[3] , 
        \u_axi4_ctrl/rfifo_wdata[4] , \u_axi4_ctrl/rfifo_wdata[5] , \u_axi4_ctrl/rfifo_wdata[6] , 
        \u_axi4_ctrl/rfifo_wdata[7] , \u_axi4_ctrl/rfifo_wdata[8] , \u_axi4_ctrl/rfifo_wdata[9] , 
        \u_axi4_ctrl/rfifo_wdata[10] , \u_axi4_ctrl/rfifo_wdata[11] , \u_axi4_ctrl/rfifo_wdata[12] , 
        \u_axi4_ctrl/rfifo_wdata[13] , \u_axi4_ctrl/rfifo_wdata[14] , \u_axi4_ctrl/rfifo_wdata[15] , 
        \u_axi4_ctrl/rfifo_wdata[16] , \u_axi4_ctrl/rfifo_wdata[17] , \u_axi4_ctrl/rfifo_wdata[18] , 
        \u_axi4_ctrl/rfifo_wdata[19] , \u_axi4_ctrl/rfifo_wdata[20] , \u_axi4_ctrl/rfifo_wdata[21] , 
        \u_axi4_ctrl/rfifo_wdata[22] , \u_axi4_ctrl/rfifo_wdata[23] , \u_axi4_ctrl/rfifo_wdata[24] , 
        \u_axi4_ctrl/rfifo_wdata[25] , \u_axi4_ctrl/rfifo_wdata[26] , \u_axi4_ctrl/rfifo_wdata[27] , 
        \u_axi4_ctrl/rfifo_wdata[28] , \u_axi4_ctrl/rfifo_wdata[29] , \u_axi4_ctrl/rfifo_wdata[30] , 
        \u_axi4_ctrl/rfifo_wdata[31] , \u_axi4_ctrl/rfifo_wdata[32] , \u_axi4_ctrl/rfifo_wdata[33] , 
        \u_axi4_ctrl/rfifo_wdata[34] , \u_axi4_ctrl/rfifo_wdata[35] , \u_axi4_ctrl/rfifo_wdata[36] , 
        \u_axi4_ctrl/rfifo_wdata[37] , \u_axi4_ctrl/rfifo_wdata[38] , \u_axi4_ctrl/rfifo_wdata[39] , 
        \u_axi4_ctrl/rfifo_wdata[40] , \u_axi4_ctrl/rfifo_wdata[41] , \u_axi4_ctrl/rfifo_wdata[42] , 
        \u_axi4_ctrl/rfifo_wdata[43] , \u_axi4_ctrl/rfifo_wdata[44] , \u_axi4_ctrl/rfifo_wdata[45] , 
        \u_axi4_ctrl/rfifo_wdata[46] , \u_axi4_ctrl/rfifo_wdata[47] , \u_axi4_ctrl/rfifo_wdata[48] , 
        \u_axi4_ctrl/rfifo_wdata[49] , \u_axi4_ctrl/rfifo_wdata[50] , \u_axi4_ctrl/rfifo_wdata[51] , 
        \u_axi4_ctrl/rfifo_wdata[52] , \u_axi4_ctrl/rfifo_wdata[53] , \u_axi4_ctrl/rfifo_wdata[54] , 
        \u_axi4_ctrl/rfifo_wdata[55] , \u_axi4_ctrl/rfifo_wdata[56] , \u_axi4_ctrl/rfifo_wdata[57] , 
        \u_axi4_ctrl/rfifo_wdata[58] , \u_axi4_ctrl/rfifo_wdata[59] , \u_axi4_ctrl/rfifo_wdata[60] , 
        \u_axi4_ctrl/rfifo_wdata[61] , \u_axi4_ctrl/rfifo_wdata[62] , \u_axi4_ctrl/rfifo_wdata[63] , 
        \u_axi4_ctrl/rfifo_wdata[64] , \u_axi4_ctrl/rfifo_wdata[65] , \u_axi4_ctrl/rfifo_wdata[66] , 
        \u_axi4_ctrl/rfifo_wdata[67] , \u_axi4_ctrl/rfifo_wdata[68] , \u_axi4_ctrl/rfifo_wdata[69] , 
        \u_axi4_ctrl/rfifo_wdata[70] , \u_axi4_ctrl/rfifo_wdata[71] , \u_axi4_ctrl/rfifo_wdata[72] , 
        \u_axi4_ctrl/rfifo_wdata[73] , \u_axi4_ctrl/rfifo_wdata[74] , \u_axi4_ctrl/rfifo_wdata[75] , 
        \u_axi4_ctrl/rfifo_wdata[76] , \u_axi4_ctrl/rfifo_wdata[77] , \u_axi4_ctrl/rfifo_wdata[78] , 
        \u_axi4_ctrl/rfifo_wdata[79] , \u_axi4_ctrl/rfifo_wdata[80] , \u_axi4_ctrl/rfifo_wdata[81] , 
        \u_axi4_ctrl/rfifo_wdata[82] , \u_axi4_ctrl/rfifo_wdata[83] , \u_axi4_ctrl/rfifo_wdata[84] , 
        \u_axi4_ctrl/rfifo_wdata[85] , \u_axi4_ctrl/rfifo_wdata[86] , \u_axi4_ctrl/rfifo_wdata[87] , 
        \u_axi4_ctrl/rfifo_wdata[88] , \u_axi4_ctrl/rfifo_wdata[89] , \u_axi4_ctrl/rfifo_wdata[90] , 
        \u_axi4_ctrl/rfifo_wdata[91] , \u_axi4_ctrl/rfifo_wdata[92] , \u_axi4_ctrl/rfifo_wdata[93] , 
        \u_axi4_ctrl/rfifo_wdata[94] , \u_axi4_ctrl/rfifo_wdata[95] , \u_axi4_ctrl/rfifo_wdata[96] , 
        \u_axi4_ctrl/rfifo_wdata[97] , \u_axi4_ctrl/rfifo_wdata[98] , \u_axi4_ctrl/rfifo_wdata[99] , 
        \u_axi4_ctrl/rfifo_wdata[100] , \u_axi4_ctrl/rfifo_wdata[101] , 
        \u_axi4_ctrl/rfifo_wdata[102] , \u_axi4_ctrl/rfifo_wdata[103] , 
        \u_axi4_ctrl/rfifo_wdata[104] , \u_axi4_ctrl/rfifo_wdata[105] , 
        \u_axi4_ctrl/rfifo_wdata[106] , \u_axi4_ctrl/rfifo_wdata[107] , 
        \u_axi4_ctrl/rfifo_wdata[108] , \u_axi4_ctrl/rfifo_wdata[109] , 
        \u_axi4_ctrl/rfifo_wdata[110] , \u_axi4_ctrl/rfifo_wdata[111] , 
        \u_axi4_ctrl/rfifo_wdata[112] , \u_axi4_ctrl/rfifo_wdata[113] , 
        \u_axi4_ctrl/rfifo_wdata[114] , \u_axi4_ctrl/rfifo_wdata[115] , 
        \u_axi4_ctrl/rfifo_wdata[116] , \u_axi4_ctrl/rfifo_wdata[117] , 
        \u_axi4_ctrl/rfifo_wdata[118] , \u_axi4_ctrl/rfifo_wdata[119] , 
        \u_axi4_ctrl/rfifo_wdata[120] , \u_axi4_ctrl/rfifo_wdata[121] , 
        \u_axi4_ctrl/rfifo_wdata[122] , \u_axi4_ctrl/rfifo_wdata[123] , 
        \u_axi4_ctrl/rfifo_wdata[124] , \u_axi4_ctrl/rfifo_wdata[125] , 
        \u_axi4_ctrl/rfifo_wdata[126] , \u_axi4_ctrl/rfifo_wdata[127] , 
        n3039, n3040, n3041, n3042, \u_lcd_driver/vcnt[0] , lcd_hs, 
        n3045, n3046, n3047, n3048, n3049, n3050, lcd_de, n3053, 
        n3054, n3055, n3056, \u_lcd_driver/r_lcd_dv , \u_lcd_driver/hcnt[0] , 
        n3060, n3061, n3062, n3063, \u_lcd_driver/vcnt[1] , \u_lcd_driver/vcnt[2] , 
        \u_lcd_driver/vcnt[3] , \u_lcd_driver/vcnt[4] , \u_lcd_driver/vcnt[5] , 
        \u_lcd_driver/vcnt[6] , \u_lcd_driver/vcnt[7] , \u_lcd_driver/vcnt[8] , 
        \u_lcd_driver/vcnt[9] , \u_lcd_driver/vcnt[10] , \u_lcd_driver/vcnt[11] , 
        n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, 
        n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, 
        n3091, n3092, \u_lcd_driver/hcnt[1] , \u_lcd_driver/hcnt[2] , 
        \u_lcd_driver/hcnt[3] , \u_lcd_driver/hcnt[4] , \u_lcd_driver/hcnt[5] , 
        \u_lcd_driver/hcnt[6] , \u_lcd_driver/hcnt[7] , \u_lcd_driver/hcnt[8] , 
        \u_lcd_driver/hcnt[9] , \u_lcd_driver/hcnt[10] , \u_lcd_driver/hcnt[11] , 
        n3203, n3204, \w_hdmi_txd0[0] , \u_rgb2dvi/enc_0/acc[0] , n3217, 
        n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, 
        n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
        n3234, n3235, n3236, n3237, \w_hdmi_txd0[1] , \w_hdmi_txd0[2] , 
        \w_hdmi_txd0[3] , \w_hdmi_txd0[4] , \w_hdmi_txd0[5] , \w_hdmi_txd0[6] , 
        \w_hdmi_txd0[7] , \w_hdmi_txd0[8] , \w_hdmi_txd0[9] , \u_rgb2dvi/enc_0/acc[1] , 
        \u_rgb2dvi/enc_0/acc[2] , \u_rgb2dvi/enc_0/acc[3] , \u_rgb2dvi/enc_0/acc[4] , 
        n3282, n3283, \w_hdmi_txd1[0] , \u_rgb2dvi/enc_1/acc[0] , n3294, 
        n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
        n3303, n3304, n3305, n3306, n3307, \w_hdmi_txd1[1] , \w_hdmi_txd1[2] , 
        \w_hdmi_txd1[3] , \w_hdmi_txd1[4] , \w_hdmi_txd1[5] , \w_hdmi_txd1[6] , 
        \w_hdmi_txd1[7] , \w_hdmi_txd1[8] , \w_hdmi_txd1[9] , n3317, 
        n3318, n3319, n3320, n3321, n3322, n3323, n3324, \u_rgb2dvi/enc_1/acc[1] , 
        \u_rgb2dvi/enc_1/acc[2] , \u_rgb2dvi/enc_1/acc[3] , \u_rgb2dvi/enc_1/acc[4] , 
        n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, 
        n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, 
        \w_hdmi_txd2[0] , n3346, n3347, n3348, n3349, \u_rgb2dvi/enc_2/acc[0] , 
        n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
        n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
        n3367, n3368, n3369, \w_hdmi_txd2[1] , \w_hdmi_txd2[2] , \w_hdmi_txd2[3] , 
        \w_hdmi_txd2[4] , \w_hdmi_txd2[5] , \w_hdmi_txd2[6] , \w_hdmi_txd2[7] , 
        \w_hdmi_txd2[9] , n3378, n3379, n3380, n3381, n3382, n3383, 
        n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, 
        n3392, n3393, \u_rgb2dvi/enc_2/acc[1] , \u_rgb2dvi/enc_2/acc[2] , 
        \u_rgb2dvi/enc_2/acc[3] , \u_rgb2dvi/enc_2/acc[4] , n3398, n3399, 
        n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, 
        n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, 
        n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, 
        n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, 
        n3432, n3433, n3434, n3436, n3437, n3438, n3439, n3440, 
        n3441, n3442, \r_hdmi_tx0_o[5] , \r_hdmi_tx0_o[6] , \r_hdmi_tx0_o[7] , 
        \r_hdmi_tx0_o[8] , \r_hdmi_tx0_o[9] , \r_hdmi_tx1_o[5] , \r_hdmi_tx1_o[6] , 
        \r_hdmi_tx1_o[7] , \r_hdmi_tx1_o[8] , \r_hdmi_tx1_o[9] , \r_hdmi_tx2_o[5] , 
        \r_hdmi_tx2_o[6] , \r_hdmi_tx2_o[7] , \r_hdmi_tx2_o[9] , \PowerOnResetCnt[1] , 
        \PowerOnResetCnt[2] , \PowerOnResetCnt[3] , \PowerOnResetCnt[4] , 
        \PowerOnResetCnt[5] , \PowerOnResetCnt[6] , \PowerOnResetCnt[7] , 
        \edb_top_inst/n1731 , \edb_top_inst/la0/la_run_trig , \edb_top_inst/la0/la_trig_pattern[0] , 
        \edb_top_inst/la0/la_run_trig_imdt , \edb_top_inst/la0/la_stop_trig , 
        \edb_top_inst/la0/la_capture_pattern[0] , \edb_top_inst/la0/la_trig_mask[0] , 
        \edb_top_inst/la0/la_num_trigger[0] , \edb_top_inst/la0/la_window_depth[0] , 
        \edb_top_inst/la0/la_soft_reset_in , \edb_top_inst/la0/address_counter[0] , 
        \edb_top_inst/la0/opcode[0] , \edb_top_inst/la0/bit_count[0] , \edb_top_inst/la0/word_count[0] , 
        \edb_top_inst/la0/data_out_shift_reg[0] , \edb_top_inst/la0/module_state[0] , 
        \edb_top_inst/la0/la_resetn_p1 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/la_resetn , \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/cap_fifo_din_cu[0] , \edb_top_inst/la0/cap_fifo_din_tu[0] , 
        \edb_top_inst/la0/internal_register_select[0] , \edb_top_inst/la0/la_trig_pos[0] , 
        \edb_top_inst/la0/la_trig_pattern[1] , \edb_top_inst/la0/la_capture_pattern[1] , 
        \edb_top_inst/la0/la_trig_mask[1] , \edb_top_inst/la0/la_trig_mask[2] , 
        \edb_top_inst/la0/la_trig_mask[3] , \edb_top_inst/la0/la_trig_mask[4] , 
        \edb_top_inst/la0/la_trig_mask[5] , \edb_top_inst/la0/la_trig_mask[6] , 
        \edb_top_inst/la0/la_trig_mask[7] , \edb_top_inst/la0/la_trig_mask[8] , 
        \edb_top_inst/la0/la_trig_mask[9] , \edb_top_inst/la0/la_trig_mask[10] , 
        \edb_top_inst/la0/la_trig_mask[11] , \edb_top_inst/la0/la_trig_mask[12] , 
        \edb_top_inst/la0/la_trig_mask[13] , \edb_top_inst/la0/la_trig_mask[14] , 
        \edb_top_inst/la0/la_trig_mask[15] , \edb_top_inst/la0/la_trig_mask[16] , 
        \edb_top_inst/la0/la_trig_mask[17] , \edb_top_inst/la0/la_trig_mask[18] , 
        \edb_top_inst/la0/la_trig_mask[19] , \edb_top_inst/la0/la_trig_mask[20] , 
        \edb_top_inst/la0/la_trig_mask[21] , \edb_top_inst/la0/la_trig_mask[22] , 
        \edb_top_inst/la0/la_trig_mask[23] , \edb_top_inst/la0/la_trig_mask[24] , 
        \edb_top_inst/la0/la_trig_mask[25] , \edb_top_inst/la0/la_trig_mask[26] , 
        \edb_top_inst/la0/la_trig_mask[27] , \edb_top_inst/la0/la_trig_mask[28] , 
        \edb_top_inst/la0/la_trig_mask[29] , \edb_top_inst/la0/la_trig_mask[30] , 
        \edb_top_inst/la0/la_trig_mask[31] , \edb_top_inst/la0/la_trig_mask[32] , 
        \edb_top_inst/la0/la_trig_mask[33] , \edb_top_inst/la0/la_trig_mask[34] , 
        \edb_top_inst/la0/la_trig_mask[35] , \edb_top_inst/la0/la_trig_mask[36] , 
        \edb_top_inst/la0/la_trig_mask[37] , \edb_top_inst/la0/la_trig_mask[38] , 
        \edb_top_inst/la0/la_trig_mask[39] , \edb_top_inst/la0/la_trig_mask[40] , 
        \edb_top_inst/la0/la_trig_mask[41] , \edb_top_inst/la0/la_trig_mask[42] , 
        \edb_top_inst/la0/la_trig_mask[43] , \edb_top_inst/la0/la_trig_mask[44] , 
        \edb_top_inst/la0/la_trig_mask[45] , \edb_top_inst/la0/la_trig_mask[46] , 
        \edb_top_inst/la0/la_trig_mask[47] , \edb_top_inst/la0/la_trig_mask[48] , 
        \edb_top_inst/la0/la_trig_mask[49] , \edb_top_inst/la0/la_trig_mask[50] , 
        \edb_top_inst/la0/la_trig_mask[51] , \edb_top_inst/la0/la_trig_mask[52] , 
        \edb_top_inst/la0/la_trig_mask[53] , \edb_top_inst/la0/la_trig_mask[54] , 
        \edb_top_inst/la0/la_trig_mask[55] , \edb_top_inst/la0/la_trig_mask[56] , 
        \edb_top_inst/la0/la_trig_mask[57] , \edb_top_inst/la0/la_trig_mask[58] , 
        \edb_top_inst/la0/la_trig_mask[59] , \edb_top_inst/la0/la_trig_mask[60] , 
        \edb_top_inst/la0/la_trig_mask[61] , \edb_top_inst/la0/la_trig_mask[62] , 
        \edb_top_inst/la0/la_trig_mask[63] , \edb_top_inst/la0/la_num_trigger[1] , 
        \edb_top_inst/la0/la_num_trigger[2] , \edb_top_inst/la0/la_num_trigger[3] , 
        \edb_top_inst/la0/la_num_trigger[4] , \edb_top_inst/la0/la_num_trigger[5] , 
        \edb_top_inst/la0/la_num_trigger[6] , \edb_top_inst/la0/la_num_trigger[7] , 
        \edb_top_inst/la0/la_num_trigger[8] , \edb_top_inst/la0/la_num_trigger[9] , 
        \edb_top_inst/la0/la_num_trigger[10] , \edb_top_inst/la0/la_num_trigger[11] , 
        \edb_top_inst/la0/la_num_trigger[12] , \edb_top_inst/la0/la_num_trigger[13] , 
        \edb_top_inst/la0/la_num_trigger[14] , \edb_top_inst/la0/la_num_trigger[15] , 
        \edb_top_inst/la0/la_num_trigger[16] , \edb_top_inst/la0/la_window_depth[1] , 
        \edb_top_inst/la0/la_window_depth[2] , \edb_top_inst/la0/la_window_depth[3] , 
        \edb_top_inst/la0/la_window_depth[4] , \edb_top_inst/la0/address_counter[1] , 
        \edb_top_inst/la0/address_counter[2] , \edb_top_inst/la0/address_counter[3] , 
        \edb_top_inst/la0/address_counter[4] , \edb_top_inst/la0/address_counter[5] , 
        \edb_top_inst/la0/address_counter[6] , \edb_top_inst/la0/address_counter[7] , 
        \edb_top_inst/la0/address_counter[8] , \edb_top_inst/la0/address_counter[9] , 
        \edb_top_inst/la0/address_counter[10] , \edb_top_inst/la0/address_counter[11] , 
        \edb_top_inst/la0/address_counter[12] , \edb_top_inst/la0/address_counter[13] , 
        \edb_top_inst/la0/address_counter[14] , \edb_top_inst/la0/address_counter[15] , 
        \edb_top_inst/la0/address_counter[16] , \edb_top_inst/la0/address_counter[17] , 
        \edb_top_inst/la0/address_counter[18] , \edb_top_inst/la0/address_counter[19] , 
        \edb_top_inst/la0/address_counter[20] , \edb_top_inst/la0/address_counter[21] , 
        \edb_top_inst/la0/address_counter[22] , \edb_top_inst/la0/address_counter[23] , 
        \edb_top_inst/la0/address_counter[24] , \edb_top_inst/la0/address_counter[25] , 
        \edb_top_inst/la0/address_counter[26] , \edb_top_inst/la0/opcode[1] , 
        \edb_top_inst/la0/opcode[2] , \edb_top_inst/la0/opcode[3] , \edb_top_inst/la0/bit_count[1] , 
        \edb_top_inst/la0/bit_count[2] , \edb_top_inst/la0/bit_count[3] , 
        \edb_top_inst/la0/bit_count[4] , \edb_top_inst/la0/bit_count[5] , 
        \edb_top_inst/la0/word_count[1] , \edb_top_inst/la0/word_count[2] , 
        \edb_top_inst/la0/word_count[3] , \edb_top_inst/la0/word_count[4] , 
        \edb_top_inst/la0/word_count[5] , \edb_top_inst/la0/word_count[6] , 
        \edb_top_inst/la0/word_count[7] , \edb_top_inst/la0/word_count[8] , 
        \edb_top_inst/la0/word_count[9] , \edb_top_inst/la0/word_count[10] , 
        \edb_top_inst/la0/word_count[11] , \edb_top_inst/la0/word_count[12] , 
        \edb_top_inst/la0/word_count[13] , \edb_top_inst/la0/word_count[14] , 
        \edb_top_inst/la0/word_count[15] , \edb_top_inst/la0/data_out_shift_reg[1] , 
        \edb_top_inst/la0/data_out_shift_reg[2] , \edb_top_inst/la0/data_out_shift_reg[3] , 
        \edb_top_inst/la0/data_out_shift_reg[4] , \edb_top_inst/la0/data_out_shift_reg[5] , 
        \edb_top_inst/la0/data_out_shift_reg[6] , \edb_top_inst/la0/data_out_shift_reg[7] , 
        \edb_top_inst/la0/data_out_shift_reg[8] , \edb_top_inst/la0/data_out_shift_reg[9] , 
        \edb_top_inst/la0/data_out_shift_reg[10] , \edb_top_inst/la0/data_out_shift_reg[11] , 
        \edb_top_inst/la0/data_out_shift_reg[12] , \edb_top_inst/la0/data_out_shift_reg[13] , 
        \edb_top_inst/la0/data_out_shift_reg[14] , \edb_top_inst/la0/data_out_shift_reg[15] , 
        \edb_top_inst/la0/data_out_shift_reg[16] , \edb_top_inst/la0/data_out_shift_reg[17] , 
        \edb_top_inst/la0/data_out_shift_reg[18] , \edb_top_inst/la0/data_out_shift_reg[19] , 
        \edb_top_inst/la0/data_out_shift_reg[20] , \edb_top_inst/la0/data_out_shift_reg[21] , 
        \edb_top_inst/la0/data_out_shift_reg[22] , \edb_top_inst/la0/data_out_shift_reg[23] , 
        \edb_top_inst/la0/data_out_shift_reg[24] , \edb_top_inst/la0/data_out_shift_reg[25] , 
        \edb_top_inst/la0/data_out_shift_reg[26] , \edb_top_inst/la0/data_out_shift_reg[27] , 
        \edb_top_inst/la0/data_out_shift_reg[28] , \edb_top_inst/la0/data_out_shift_reg[29] , 
        \edb_top_inst/la0/data_out_shift_reg[30] , \edb_top_inst/la0/data_out_shift_reg[31] , 
        \edb_top_inst/la0/data_out_shift_reg[32] , \edb_top_inst/la0/data_out_shift_reg[33] , 
        \edb_top_inst/la0/data_out_shift_reg[34] , \edb_top_inst/la0/data_out_shift_reg[35] , 
        \edb_top_inst/la0/data_out_shift_reg[36] , \edb_top_inst/la0/data_out_shift_reg[37] , 
        \edb_top_inst/la0/data_out_shift_reg[38] , \edb_top_inst/la0/data_out_shift_reg[39] , 
        \edb_top_inst/la0/data_out_shift_reg[40] , \edb_top_inst/la0/data_out_shift_reg[41] , 
        \edb_top_inst/la0/data_out_shift_reg[42] , \edb_top_inst/la0/data_out_shift_reg[43] , 
        \edb_top_inst/la0/data_out_shift_reg[44] , \edb_top_inst/la0/data_out_shift_reg[45] , 
        \edb_top_inst/la0/data_out_shift_reg[46] , \edb_top_inst/la0/data_out_shift_reg[47] , 
        \edb_top_inst/la0/data_out_shift_reg[48] , \edb_top_inst/la0/data_out_shift_reg[49] , 
        \edb_top_inst/la0/data_out_shift_reg[50] , \edb_top_inst/la0/data_out_shift_reg[51] , 
        \edb_top_inst/la0/data_out_shift_reg[52] , \edb_top_inst/la0/data_out_shift_reg[53] , 
        \edb_top_inst/la0/data_out_shift_reg[54] , \edb_top_inst/la0/data_out_shift_reg[55] , 
        \edb_top_inst/la0/data_out_shift_reg[56] , \edb_top_inst/la0/data_out_shift_reg[57] , 
        \edb_top_inst/la0/data_out_shift_reg[58] , \edb_top_inst/la0/data_out_shift_reg[59] , 
        \edb_top_inst/la0/data_out_shift_reg[60] , \edb_top_inst/la0/data_out_shift_reg[61] , 
        \edb_top_inst/la0/data_out_shift_reg[62] , \edb_top_inst/la0/data_out_shift_reg[63] , 
        \edb_top_inst/la0/module_state[1] , \edb_top_inst/la0/module_state[2] , 
        \edb_top_inst/la0/module_state[3] , \edb_top_inst/la0/crc_data_out[0] , 
        \edb_top_inst/la0/crc_data_out[1] , \edb_top_inst/la0/crc_data_out[2] , 
        \edb_top_inst/la0/crc_data_out[3] , \edb_top_inst/la0/crc_data_out[4] , 
        \edb_top_inst/la0/crc_data_out[5] , \edb_top_inst/la0/crc_data_out[6] , 
        \edb_top_inst/la0/crc_data_out[7] , \edb_top_inst/la0/crc_data_out[8] , 
        \edb_top_inst/la0/crc_data_out[9] , \edb_top_inst/la0/crc_data_out[10] , 
        \edb_top_inst/la0/crc_data_out[11] , \edb_top_inst/la0/crc_data_out[12] , 
        \edb_top_inst/la0/crc_data_out[13] , \edb_top_inst/la0/crc_data_out[14] , 
        \edb_top_inst/la0/crc_data_out[15] , \edb_top_inst/la0/crc_data_out[16] , 
        \edb_top_inst/la0/crc_data_out[17] , \edb_top_inst/la0/crc_data_out[18] , 
        \edb_top_inst/la0/crc_data_out[19] , \edb_top_inst/la0/crc_data_out[20] , 
        \edb_top_inst/la0/crc_data_out[21] , \edb_top_inst/la0/crc_data_out[22] , 
        \edb_top_inst/la0/crc_data_out[23] , \edb_top_inst/la0/crc_data_out[24] , 
        \edb_top_inst/la0/crc_data_out[25] , \edb_top_inst/la0/crc_data_out[26] , 
        \edb_top_inst/la0/crc_data_out[27] , \edb_top_inst/la0/crc_data_out[28] , 
        \edb_top_inst/la0/crc_data_out[29] , \edb_top_inst/la0/crc_data_out[30] , 
        \edb_top_inst/la0/crc_data_out[31] , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/tu_trigger , \edb_top_inst/la0/cap_fifo_din_cu[1] , 
        \edb_top_inst/la0/cap_fifo_din_cu[2] , \edb_top_inst/la0/cap_fifo_din_cu[3] , 
        \edb_top_inst/la0/cap_fifo_din_cu[4] , \edb_top_inst/la0/cap_fifo_din_cu[5] , 
        \edb_top_inst/la0/cap_fifo_din_cu[6] , \edb_top_inst/la0/cap_fifo_din_cu[7] , 
        \edb_top_inst/la0/cap_fifo_din_cu[8] , \edb_top_inst/la0/cap_fifo_din_cu[9] , 
        \edb_top_inst/la0/cap_fifo_din_tu[1] , \edb_top_inst/la0/cap_fifo_din_tu[2] , 
        \edb_top_inst/la0/cap_fifo_din_tu[3] , \edb_top_inst/la0/cap_fifo_din_tu[4] , 
        \edb_top_inst/la0/cap_fifo_din_tu[5] , \edb_top_inst/la0/cap_fifo_din_tu[6] , 
        \edb_top_inst/la0/cap_fifo_din_tu[7] , \edb_top_inst/la0/cap_fifo_din_tu[8] , 
        \edb_top_inst/la0/cap_fifo_din_tu[9] , \edb_top_inst/la0/la_biu_inst/curr_state[0] , 
        \edb_top_inst/la0/la_biu_inst/run_trig_p2 , \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 , 
        \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 , \edb_top_inst/la0/la_biu_inst/str_sync , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff1 , \edb_top_inst/la0/la_biu_inst/str_sync_wbff2 , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q , \edb_top_inst/la0/la_biu_inst/rdy_sync , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q , \edb_top_inst/la0/data_from_biu[0] , 
        \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] , \edb_top_inst/la0/la_biu_inst/curr_state[3] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[2] , \edb_top_inst/la0/la_biu_inst/curr_state[1] , 
        \edb_top_inst/la0/biu_ready , \edb_top_inst/la0/la_biu_inst/addr_reg[15] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[16] , \edb_top_inst/la0/la_biu_inst/addr_reg[17] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[18] , \edb_top_inst/la0/la_biu_inst/addr_reg[19] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[20] , \edb_top_inst/la0/la_biu_inst/addr_reg[21] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[22] , \edb_top_inst/la0/la_biu_inst/addr_reg[23] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[24] , \edb_top_inst/la0/la_biu_inst/addr_reg[25] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[26] , \edb_top_inst/la0/data_from_biu[1] , 
        \edb_top_inst/la0/data_from_biu[2] , \edb_top_inst/la0/data_from_biu[3] , 
        \edb_top_inst/la0/data_from_biu[4] , \edb_top_inst/la0/data_from_biu[5] , 
        \edb_top_inst/la0/data_from_biu[6] , \edb_top_inst/la0/data_from_biu[7] , 
        \edb_top_inst/la0/data_from_biu[8] , \edb_top_inst/la0/data_from_biu[9] , 
        \edb_top_inst/la0/data_from_biu[10] , \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] , 
        \edb_top_inst/la0/la_sample_cnt[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[0] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] , 
        \edb_top_inst/la0/la_sample_cnt[1] , \edb_top_inst/la0/la_sample_cnt[2] , 
        \edb_top_inst/la0/la_sample_cnt[3] , \edb_top_inst/la0/la_sample_cnt[4] , 
        \edb_top_inst/la0/la_sample_cnt[5] , \edb_top_inst/la0/la_sample_cnt[6] , 
        \edb_top_inst/la0/la_sample_cnt[7] , \edb_top_inst/la0/la_sample_cnt[8] , 
        \edb_top_inst/la0/la_sample_cnt[9] , \edb_top_inst/la0/la_sample_cnt[10] , 
        \edb_top_inst/la0/la_sample_cnt[11] , \edb_top_inst/la0/la_sample_cnt[12] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[1] , \edb_top_inst/la0/la_biu_inst/fifo_counter[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[3] , \edb_top_inst/la0/la_biu_inst/fifo_counter[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[5] , \edb_top_inst/la0/la_biu_inst/fifo_counter[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[7] , \edb_top_inst/la0/la_biu_inst/fifo_counter[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[9] , \edb_top_inst/la0/la_biu_inst/fifo_counter[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[11] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] , 
        \edb_top_inst/la0/internal_register_select[1] , \edb_top_inst/la0/internal_register_select[2] , 
        \edb_top_inst/la0/internal_register_select[3] , \edb_top_inst/la0/internal_register_select[4] , 
        \edb_top_inst/la0/internal_register_select[5] , \edb_top_inst/la0/internal_register_select[6] , 
        \edb_top_inst/la0/internal_register_select[7] , \edb_top_inst/la0/internal_register_select[8] , 
        \edb_top_inst/la0/internal_register_select[9] , \edb_top_inst/la0/internal_register_select[10] , 
        \edb_top_inst/la0/internal_register_select[11] , \edb_top_inst/la0/internal_register_select[12] , 
        \edb_top_inst/la0/la_trig_pos[1] , \edb_top_inst/la0/la_trig_pos[2] , 
        \edb_top_inst/la0/la_trig_pos[3] , \edb_top_inst/la0/la_trig_pos[4] , 
        \edb_top_inst/la0/la_trig_pos[5] , \edb_top_inst/la0/la_trig_pos[6] , 
        \edb_top_inst/la0/la_trig_pos[7] , \edb_top_inst/la0/la_trig_pos[8] , 
        \edb_top_inst/la0/la_trig_pos[9] , \edb_top_inst/la0/la_trig_pos[10] , 
        \edb_top_inst/la0/la_trig_pos[11] , \edb_top_inst/la0/la_trig_pos[12] , 
        \edb_top_inst/la0/la_trig_pos[13] , \edb_top_inst/la0/la_trig_pos[14] , 
        \edb_top_inst/la0/la_trig_pos[15] , \edb_top_inst/la0/la_trig_pos[16] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[0] , \edb_top_inst/debug_hub_inst/module_id_reg[1] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[2] , \edb_top_inst/debug_hub_inst/module_id_reg[3] , 
        \edb_top_inst/n35 , \edb_top_inst/n37 , \edb_top_inst/n298 , \edb_top_inst/n427 , 
        \edb_top_inst/n429 , \edb_top_inst/n433 , \edb_top_inst/n435 , 
        \edb_top_inst/n1732 , \edb_top_inst/n1733 , \edb_top_inst/n1734 , 
        \edb_top_inst/n1735 , \edb_top_inst/n1736 , \edb_top_inst/n1737 , 
        \edb_top_inst/n1738 , \edb_top_inst/n1739 , \edb_top_inst/n1740 , 
        \edb_top_inst/n1741 , \edb_top_inst/n1742 , \edb_top_inst/n1743 , 
        \edb_top_inst/n1744 , \edb_top_inst/n1745 , \edb_top_inst/n1746 , 
        \edb_top_inst/n1747 , \edb_top_inst/n1748 , \edb_top_inst/n1749 , 
        \edb_top_inst/n1750 , \edb_top_inst/n1751 , \edb_top_inst/n1752 , 
        \edb_top_inst/n1753 , \edb_top_inst/n1754 , \edb_top_inst/n1755 , 
        \edb_top_inst/n1756 , \edb_top_inst/n1757 , \edb_top_inst/n1758 , 
        \edb_top_inst/n1759 , \edb_top_inst/n1760 , \edb_top_inst/n1761 , 
        \edb_top_inst/n1762 , \edb_top_inst/n1763 , \edb_top_inst/n1764 , 
        \edb_top_inst/n1765 , \edb_top_inst/n1766 , \edb_top_inst/n1767 , 
        \edb_top_inst/n1768 , \edb_top_inst/n1769 , \edb_top_inst/n1770 , 
        \edb_top_inst/n1771 , \edb_top_inst/n1772 , \edb_top_inst/n1773 , 
        \edb_top_inst/n1774 , \edb_top_inst/n1775 , \edb_top_inst/n1776 , 
        \edb_top_inst/n1777 , \edb_top_inst/n1778 , \edb_top_inst/n1779 , 
        \edb_top_inst/n1780 , \edb_top_inst/n1781 , \edb_top_inst/n1782 , 
        \edb_top_inst/n1783 , \edb_top_inst/n1784 , \edb_top_inst/n1785 , 
        \edb_top_inst/n1786 , \edb_top_inst/n1787 , \edb_top_inst/n1788 , 
        \edb_top_inst/n1789 , \edb_top_inst/n1790 , \edb_top_inst/n1708 , 
        \edb_top_inst/n1705 , \edb_top_inst/n1791 , \edb_top_inst/n1792 , 
        \edb_top_inst/n1793 , \edb_top_inst/n1794 , \edb_top_inst/n1795 , 
        \edb_top_inst/n1796 , \edb_top_inst/n1797 , \edb_top_inst/n1798 , 
        \edb_top_inst/n1799 , \edb_top_inst/n1800 , \edb_top_inst/n1801 , 
        \edb_top_inst/n969 , \edb_top_inst/n1802 , \edb_top_inst/n1803 , 
        \edb_top_inst/n1804 , \edb_top_inst/n1805 , \edb_top_inst/n1806 , 
        \edb_top_inst/n1807 , \edb_top_inst/n1808 , \edb_top_inst/n1809 , 
        \edb_top_inst/n1810 , \edb_top_inst/n1811 , \edb_top_inst/n1812 , 
        \edb_top_inst/n1813 , \edb_top_inst/n1814 , \edb_top_inst/n1815 , 
        \edb_top_inst/n1816 , \edb_top_inst/n1817 , \edb_top_inst/n1818 , 
        \edb_top_inst/n1819 , \edb_top_inst/n1820 , \edb_top_inst/n1821 , 
        \edb_top_inst/n1822 , \edb_top_inst/n1823 , \edb_top_inst/n1824 , 
        \edb_top_inst/n1825 , \edb_top_inst/n1826 , \edb_top_inst/n1827 , 
        \edb_top_inst/n1828 , \edb_top_inst/n1829 , \edb_top_inst/n1830 , 
        \edb_top_inst/n1831 , \edb_top_inst/n1832 , \edb_top_inst/n1833 , 
        \edb_top_inst/n1834 , \edb_top_inst/n1835 , \edb_top_inst/n1836 , 
        \edb_top_inst/n1837 , \edb_top_inst/n1838 , \edb_top_inst/n1839 , 
        \edb_top_inst/n1840 , \edb_top_inst/n1841 , \edb_top_inst/n1842 , 
        \edb_top_inst/n1843 , \edb_top_inst/n1844 , \edb_top_inst/n1845 , 
        \edb_top_inst/n1851 , \edb_top_inst/n1852 , \edb_top_inst/n1853 , 
        \edb_top_inst/n1854 , \edb_top_inst/n1855 , \edb_top_inst/n1856 , 
        \edb_top_inst/n1857 , \edb_top_inst/n1858 , \edb_top_inst/n1859 , 
        \edb_top_inst/n1860 , \edb_top_inst/n1861 , \edb_top_inst/n1862 , 
        \edb_top_inst/n1863 , \edb_top_inst/n1864 , \edb_top_inst/n1865 , 
        \edb_top_inst/n1866 , \edb_top_inst/n1867 , \edb_top_inst/n1868 , 
        \edb_top_inst/n1869 , \edb_top_inst/n1870 , \edb_top_inst/n1871 , 
        \edb_top_inst/n1872 , \edb_top_inst/n1873 , \edb_top_inst/n1874 , 
        \edb_top_inst/n1875 , \edb_top_inst/n1876 , \edb_top_inst/n1877 , 
        \edb_top_inst/n1878 , \edb_top_inst/n1879 , \edb_top_inst/n1880 , 
        \edb_top_inst/n1881 , \edb_top_inst/n1882 , \edb_top_inst/n1883 , 
        \edb_top_inst/n1884 , \edb_top_inst/n1885 , \edb_top_inst/n1886 , 
        \edb_top_inst/n1887 , \edb_top_inst/n1888 , \edb_top_inst/n1889 , 
        \edb_top_inst/n1890 , \edb_top_inst/n1891 , \edb_top_inst/n1892 , 
        \edb_top_inst/n1893 , \edb_top_inst/n1894 , \edb_top_inst/n1895 , 
        \edb_top_inst/n1896 , \edb_top_inst/n1897 , \edb_top_inst/n1898 , 
        \edb_top_inst/n1899 , \edb_top_inst/n1900 , \edb_top_inst/n1901 , 
        \edb_top_inst/n1902 , \edb_top_inst/n1903 , \edb_top_inst/n1904 , 
        \edb_top_inst/n1905 , \edb_top_inst/n1906 , \edb_top_inst/n1907 , 
        \edb_top_inst/n1908 , \edb_top_inst/n1909 , \edb_top_inst/n1910 , 
        \edb_top_inst/n1911 , \edb_top_inst/n1912 , \edb_top_inst/n1913 , 
        \edb_top_inst/n1914 , \edb_top_inst/n1915 , \edb_top_inst/n1916 , 
        \edb_top_inst/n1917 , \edb_top_inst/n1918 , \edb_top_inst/n1919 , 
        \edb_top_inst/n1920 , \edb_top_inst/n1921 , \edb_top_inst/n1922 , 
        \edb_top_inst/n1923 , \edb_top_inst/n1924 , \edb_top_inst/n1925 , 
        \edb_top_inst/n1926 , \edb_top_inst/n1927 , \edb_top_inst/n1928 , 
        \edb_top_inst/n1929 , \edb_top_inst/n1930 , \edb_top_inst/n1931 , 
        \edb_top_inst/n1932 , \edb_top_inst/n1933 , \edb_top_inst/n1934 , 
        \edb_top_inst/n1935 , \edb_top_inst/n1936 , \edb_top_inst/n1937 , 
        \edb_top_inst/n1938 , \edb_top_inst/n1939 , \edb_top_inst/n1940 , 
        \edb_top_inst/n1941 , \edb_top_inst/n1942 , \edb_top_inst/n1943 , 
        \edb_top_inst/n1944 , \edb_top_inst/n1945 , \edb_top_inst/n1946 , 
        \edb_top_inst/n1947 , \edb_top_inst/n1948 , \edb_top_inst/n1949 , 
        \edb_top_inst/n1950 , \edb_top_inst/n1951 , \edb_top_inst/n1952 , 
        \edb_top_inst/n1953 , \edb_top_inst/n1954 , \edb_top_inst/n1955 , 
        \edb_top_inst/n1956 , \edb_top_inst/n1957 , \edb_top_inst/n1958 , 
        \edb_top_inst/n1959 , \edb_top_inst/n1960 , \edb_top_inst/n1961 , 
        \edb_top_inst/n1962 , \edb_top_inst/n1963 , \edb_top_inst/n1964 , 
        \edb_top_inst/n1965 , \edb_top_inst/n1966 , \edb_top_inst/n1967 , 
        \edb_top_inst/n1968 , \edb_top_inst/n1969 , \edb_top_inst/n1970 , 
        \edb_top_inst/n1971 , \edb_top_inst/n1972 , \edb_top_inst/n1973 , 
        \edb_top_inst/n1974 , \edb_top_inst/n1975 , \edb_top_inst/n1976 , 
        \edb_top_inst/n1977 , \edb_top_inst/n1978 , \edb_top_inst/n1979 , 
        \edb_top_inst/n1980 , \edb_top_inst/n1981 , \edb_top_inst/n1982 , 
        \edb_top_inst/n1983 , \edb_top_inst/n1984 , \edb_top_inst/n1985 , 
        \edb_top_inst/n1986 , \edb_top_inst/n1987 , \edb_top_inst/n1988 , 
        \edb_top_inst/n1989 , \edb_top_inst/n1990 , \edb_top_inst/n1991 , 
        \edb_top_inst/n1992 , \edb_top_inst/n1993 , \edb_top_inst/n1994 , 
        \edb_top_inst/n1995 , \edb_top_inst/n1996 , \edb_top_inst/n1997 , 
        \edb_top_inst/n1998 , \edb_top_inst/n1999 , \edb_top_inst/n2000 , 
        \edb_top_inst/n2001 , \edb_top_inst/n2002 , \edb_top_inst/n2003 , 
        \edb_top_inst/n2004 , \edb_top_inst/n2005 , \edb_top_inst/n2006 , 
        \edb_top_inst/n2007 , \edb_top_inst/n2008 , \edb_top_inst/n2009 , 
        \edb_top_inst/n2010 , \edb_top_inst/n2011 , \edb_top_inst/n2012 , 
        \edb_top_inst/n2013 , \edb_top_inst/n2014 , \edb_top_inst/n2015 , 
        \edb_top_inst/n2016 , \edb_top_inst/n2017 , \edb_top_inst/n2018 , 
        \edb_top_inst/n2019 , \edb_top_inst/n2020 , \edb_top_inst/n2021 , 
        \edb_top_inst/n2022 , \edb_top_inst/n2023 , \edb_top_inst/n2024 , 
        \edb_top_inst/n2025 , \edb_top_inst/n2026 , \edb_top_inst/n2027 , 
        \edb_top_inst/n2028 , \edb_top_inst/n2029 , \edb_top_inst/n2030 , 
        \edb_top_inst/n2031 , \edb_top_inst/n2032 , \edb_top_inst/n2033 , 
        \edb_top_inst/n2034 , \edb_top_inst/n2035 , \edb_top_inst/n2036 , 
        \edb_top_inst/n2037 , \edb_top_inst/n2038 , \edb_top_inst/n2039 , 
        \edb_top_inst/n2040 , \edb_top_inst/n2041 , \edb_top_inst/n2042 , 
        \edb_top_inst/n2043 , \edb_top_inst/n2044 , \edb_top_inst/n2045 , 
        \edb_top_inst/n2046 , \edb_top_inst/n2047 , \edb_top_inst/n2048 , 
        \edb_top_inst/n2049 , \edb_top_inst/n2050 , \edb_top_inst/n2051 , 
        \edb_top_inst/n2052 , \edb_top_inst/n2053 , \edb_top_inst/n2054 , 
        \edb_top_inst/n2055 , \edb_top_inst/n2056 , \edb_top_inst/n2057 , 
        \edb_top_inst/n2058 , \edb_top_inst/n2059 , \edb_top_inst/n2060 , 
        \edb_top_inst/n2061 , \edb_top_inst/n2062 , \edb_top_inst/n2063 , 
        \edb_top_inst/n2064 , \edb_top_inst/n2065 , \edb_top_inst/n2066 , 
        \edb_top_inst/n2067 , \edb_top_inst/n2068 , \edb_top_inst/n2069 , 
        \edb_top_inst/n2070 , \edb_top_inst/n2071 , \edb_top_inst/n2072 , 
        \edb_top_inst/n2073 , \edb_top_inst/n2074 , \edb_top_inst/n2075 , 
        \edb_top_inst/n2076 , \edb_top_inst/n2077 , \edb_top_inst/n2078 , 
        \edb_top_inst/n2079 , \edb_top_inst/n2080 , \edb_top_inst/n2081 , 
        \edb_top_inst/n2082 , \edb_top_inst/n2083 , \edb_top_inst/n2084 , 
        \edb_top_inst/n2085 , \edb_top_inst/n2086 , \edb_top_inst/n2087 , 
        \edb_top_inst/n2088 , \edb_top_inst/n2089 , \edb_top_inst/n2090 , 
        \edb_top_inst/n2091 , \edb_top_inst/n2092 , \edb_top_inst/n2093 , 
        \edb_top_inst/n2094 , \edb_top_inst/n2095 , \edb_top_inst/n2096 , 
        \edb_top_inst/n2097 , \edb_top_inst/n2098 , \edb_top_inst/n2099 , 
        \edb_top_inst/n2100 , \edb_top_inst/n2101 , \edb_top_inst/n2102 , 
        \edb_top_inst/n2103 , \edb_top_inst/n2104 , \edb_top_inst/n2105 , 
        \edb_top_inst/n2106 , \edb_top_inst/n2107 , \edb_top_inst/n2108 , 
        \edb_top_inst/n2109 , \edb_top_inst/n2110 , \edb_top_inst/n2111 , 
        \edb_top_inst/n2112 , \edb_top_inst/n2113 , \edb_top_inst/n2114 , 
        \edb_top_inst/n2115 , \edb_top_inst/n2116 , \edb_top_inst/n2117 , 
        \edb_top_inst/n2118 , \edb_top_inst/n2119 , \edb_top_inst/n2120 , 
        \edb_top_inst/n2121 , \edb_top_inst/n2122 , \edb_top_inst/n2123 , 
        \edb_top_inst/n2124 , \edb_top_inst/n2125 , \edb_top_inst/n2126 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , \edb_top_inst/n2127 , 
        \edb_top_inst/n2128 , \edb_top_inst/n2129 , \edb_top_inst/n2130 , 
        \edb_top_inst/n2131 , \edb_top_inst/n2132 , \edb_top_inst/n2133 , 
        \edb_top_inst/n2134 , \edb_top_inst/n2135 , \edb_top_inst/n2136 , 
        \edb_top_inst/n2137 , \edb_top_inst/n2138 , \edb_top_inst/n2139 , 
        \edb_top_inst/n2140 , \edb_top_inst/n2141 , \edb_top_inst/n2142 , 
        \edb_top_inst/n2143 , \edb_top_inst/n2144 , \edb_top_inst/n2145 , 
        \edb_top_inst/n2146 , \edb_top_inst/n2147 , \edb_top_inst/n2148 , 
        \edb_top_inst/n2149 , \edb_top_inst/n2150 , \edb_top_inst/n2151 , 
        \edb_top_inst/n2152 , \edb_top_inst/n2153 , \edb_top_inst/n2154 , 
        \edb_top_inst/n2155 , \edb_top_inst/n2156 , \edb_top_inst/n2157 , 
        \edb_top_inst/n2158 , \edb_top_inst/n2159 , \edb_top_inst/n2160 , 
        \edb_top_inst/n2161 , \edb_top_inst/n2162 , \edb_top_inst/n2163 , 
        \edb_top_inst/n2164 , \edb_top_inst/n2165 , \edb_top_inst/n2166 , 
        \edb_top_inst/n2167 , \edb_top_inst/n2168 , \edb_top_inst/n2169 , 
        \edb_top_inst/n2170 , \edb_top_inst/n2171 , \edb_top_inst/n2172 , 
        \edb_top_inst/n2173 , \edb_top_inst/n1711 , n4984, n4985, n4986, 
        n4987, n4988, n4989, n4990, n4991, \reduce_nand_9/n7 , DdrInitDone, 
        \Axi0ResetReg[2] , \U0_DDR_Reset/u_ddr_reset_sequencer/n15 , \U0_DDR_Reset/u_ddr_reset_sequencer/equal_21/n3 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] , \U0_DDR_Reset/u_ddr_reset_sequencer/n92 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n91 , \u_i2c_timing_ctrl_16reg_16bit/n137 , 
        \u_i2c_timing_ctrl_16reg_16bit/next_state[0] , \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en , 
        \u_i2c_timing_ctrl_16reg_16bit/n138 , \u_i2c_timing_ctrl_16reg_16bit/n139 , 
        \u_i2c_timing_ctrl_16reg_16bit/n140 , \u_i2c_timing_ctrl_16reg_16bit/n205 , 
        \u_i2c_timing_ctrl_16reg_16bit/n846 , \u_i2c_timing_ctrl_16reg_16bit/n500 , 
        ceg_net552, \u_i2c_timing_ctrl_16reg_16bit/n509 , ceg_net664, 
        \u_i2c_timing_ctrl_16reg_16bit/n567 , \u_i2c_timing_ctrl_16reg_16bit/n570 , 
        \u_i2c_timing_ctrl_16reg_16bit/n573 , \u_i2c_timing_ctrl_16reg_16bit/n576 , 
        \u_i2c_timing_ctrl_16reg_16bit/n579 , \u_i2c_timing_ctrl_16reg_16bit/n581 , 
        \u_i2c_timing_ctrl_16reg_16bit/n7 , \u_i2c_timing_ctrl_16reg_16bit/n495 , 
        ceg_net632, \u_i2c_timing_ctrl_16reg_16bit/n136 , \u_i2c_timing_ctrl_16reg_16bit/n135 , 
        \u_i2c_timing_ctrl_16reg_16bit/n134 , \u_i2c_timing_ctrl_16reg_16bit/n133 , 
        \u_i2c_timing_ctrl_16reg_16bit/n132 , \u_i2c_timing_ctrl_16reg_16bit/n131 , 
        \u_i2c_timing_ctrl_16reg_16bit/n130 , \u_i2c_timing_ctrl_16reg_16bit/n129 , 
        \u_i2c_timing_ctrl_16reg_16bit/n128 , \u_i2c_timing_ctrl_16reg_16bit/n127 , 
        \u_i2c_timing_ctrl_16reg_16bit/n126 , \u_i2c_timing_ctrl_16reg_16bit/n125 , 
        \u_i2c_timing_ctrl_16reg_16bit/n124 , \u_i2c_timing_ctrl_16reg_16bit/n123 , 
        \u_i2c_timing_ctrl_16reg_16bit/n122 , \u_i2c_timing_ctrl_16reg_16bit/next_state[1] , 
        \u_i2c_timing_ctrl_16reg_16bit/next_state[2] , \u_i2c_timing_ctrl_16reg_16bit/next_state[3] , 
        \u_i2c_timing_ctrl_16reg_16bit/next_state[4] , \u_i2c_timing_ctrl_16reg_16bit/n204 , 
        \u_i2c_timing_ctrl_16reg_16bit/n203 , \u_i2c_timing_ctrl_16reg_16bit/n202 , 
        \u_i2c_timing_ctrl_16reg_16bit/n201 , \u_i2c_timing_ctrl_16reg_16bit/n200 , 
        \u_i2c_timing_ctrl_16reg_16bit/n199 , \u_i2c_timing_ctrl_16reg_16bit/n198 , 
        \u_i2c_timing_ctrl_16reg_16bit/n499 , \u_i2c_timing_ctrl_16reg_16bit/n498 , 
        \u_i2c_timing_ctrl_16reg_16bit/n497 , \u_i2c_timing_ctrl_16reg_16bit/n508 , 
        \u_i2c_timing_ctrl_16reg_16bit/n507 , \u_i2c_timing_ctrl_16reg_16bit/n506 , 
        \u_i2c_timing_ctrl_16reg_16bit/n505 , \u_i2c_timing_ctrl_16reg_16bit/n504 , 
        \u_i2c_timing_ctrl_16reg_16bit/n503 , \u_i2c_timing_ctrl_16reg_16bit/n502 , 
        n5371, n5374, n5377, n5380, n5385, n5388, n5391, n5394, 
        n5403, n5410, n5413, n5416, n5417, n5420, n5422, n5425, 
        n5428, n5431, \u_CMOS_Capture_RAW_Gray/n127 , ceg_net126, \u_CMOS_Capture_RAW_Gray/n160 , 
        ceg_net154, \u_CMOS_Capture_RAW_Gray/n171 , \u_CMOS_Capture_RAW_Gray/n126 , 
        \u_CMOS_Capture_RAW_Gray/n125 , \u_CMOS_Capture_RAW_Gray/n124 , 
        \u_CMOS_Capture_RAW_Gray/n123 , \u_CMOS_Capture_RAW_Gray/n122 , 
        \u_CMOS_Capture_RAW_Gray/n121 , \u_CMOS_Capture_RAW_Gray/n120 , 
        \u_CMOS_Capture_RAW_Gray/n119 , \u_CMOS_Capture_RAW_Gray/n118 , 
        \u_CMOS_Capture_RAW_Gray/n117 , \u_CMOS_Capture_RAW_Gray/n116 , 
        \u_CMOS_Capture_RAW_Gray/n159 , n5623, n5626, cmos_frame_href, 
        n5660, \u_sensor_frame_count/cmos_fps_cnt[1] , \u_sensor_frame_count/n141 , 
        ceg_net200, n2090, \cmos_frame_Gray[0] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 , 
        \u_sensor_frame_count/n110 , \u_sensor_frame_count/n75 , \u_sensor_frame_count/n74 , 
        \u_sensor_frame_count/n73 , \u_sensor_frame_count/n72 , \u_sensor_frame_count/n71 , 
        \u_sensor_frame_count/n70 , \u_sensor_frame_count/n69 , \u_sensor_frame_count/n68 , 
        \u_sensor_frame_count/n67 , \u_sensor_frame_count/n66 , \u_sensor_frame_count/n65 , 
        \u_sensor_frame_count/n64 , \u_sensor_frame_count/n63 , \u_sensor_frame_count/n62 , 
        \u_sensor_frame_count/n61 , \u_sensor_frame_count/n60 , \u_sensor_frame_count/n59 , 
        \u_sensor_frame_count/n58 , \u_sensor_frame_count/n57 , \u_sensor_frame_count/n56 , 
        \u_sensor_frame_count/n55 , \u_sensor_frame_count/n54 , \u_sensor_frame_count/n53 , 
        \u_sensor_frame_count/n52 , \u_sensor_frame_count/n51 , \u_sensor_frame_count/n50 , 
        \u_sensor_frame_count/n49 , \u_sensor_frame_count/n48 , n5723, 
        \u_sensor_frame_count/n140 , \u_sensor_frame_count/n139 , \u_sensor_frame_count/n138 , 
        \u_sensor_frame_count/n137 , \u_sensor_frame_count/n136 , \u_sensor_frame_count/n135 , 
        \u_sensor_frame_count/n134 , \u_sensor_frame_count/n133 , n5734, 
        n5737, n5740, \u_afifo_buf/u_efx_fifo_top/raddr[12] , \u_afifo_buf/u_efx_fifo_top/rd_en_int , 
        n2104, \cmos_frame_Gray[2] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 , 
        \cmos_frame_Gray[1] , \cmos_frame_Gray[3] , \cmos_frame_Gray[4] , 
        \cmos_frame_Gray[5] , \cmos_frame_Gray[6] , \cmos_frame_Gray[7] , 
        \u_afifo_buf/u_efx_fifo_top/wr_en_int , ceg_net219, n5807, \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[13] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[12] , 
        ceg_net226, \u_scaler_gray/n150 , ceg_net229, tvalid_o, \u_scaler_gray/u0_data_stream_ctr/w_image_tlast , 
        \u_scaler_gray/u0_data_stream_ctr/n1703 , n197, \u_scaler_gray/u0_data_stream_ctr/n1704 , 
        \u_scaler_gray/u0_data_stream_ctr/n432 , \u_scaler_gray/u0_data_stream_ctr/n2157 , 
        ceg_net526, \u_scaler_gray/u0_data_stream_ctr/equal_59/n5 , \u_scaler_gray/u0_data_stream_ctr/n1712 , 
        \u_scaler_gray/u0_data_stream_ctr/r_image_tlast , \u_scaler_gray/u0_data_stream_ctr/n1713 , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
        \tdata_i[6] , \u_scaler_gray/u0_data_stream_ctr/n903 , \tdata_i[1] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
        \u_scaler_gray/u0_data_stream_ctr/n1702 , \u_scaler_gray/u0_data_stream_ctr/n431 , 
        \u_scaler_gray/u0_data_stream_ctr/n430 , \u_scaler_gray/u0_data_stream_ctr/n2080 , 
        \u_scaler_gray/u0_data_stream_ctr/n1162 , \u_scaler_gray/u0_data_stream_ctr/n1161 , 
        \u_scaler_gray/u0_data_stream_ctr/n1160 , \u_scaler_gray/u0_data_stream_ctr/n1159 , 
        \u_scaler_gray/u0_data_stream_ctr/n885 , \u_scaler_gray/u0_data_stream_ctr/n884 , 
        \u_scaler_gray/u0_data_stream_ctr/n883 , \u_scaler_gray/u0_data_stream_ctr/n882 , 
        \u_scaler_gray/u0_data_stream_ctr/n881 , \u_scaler_gray/u0_data_stream_ctr/n880 , 
        \u_scaler_gray/u0_data_stream_ctr/n879 , \u_scaler_gray/u0_data_stream_ctr/n1179 , 
        \u_scaler_gray/u0_data_stream_ctr/n1178 , \u_scaler_gray/u0_data_stream_ctr/n1177 , 
        \u_scaler_gray/u0_data_stream_ctr/n1176 , \u_scaler_gray/u0_data_stream_ctr/n1195 , 
        \u_scaler_gray/u0_data_stream_ctr/n1194 , \u_scaler_gray/u0_data_stream_ctr/n1193 , 
        \u_scaler_gray/u0_data_stream_ctr/n1212 , \u_scaler_gray/u0_data_stream_ctr/n1211 , 
        \u_scaler_gray/u0_data_stream_ctr/n1210 , \tdata_i[5] , \tdata_i[7] , 
        \tdata_i[4] , \tdata_i[2] , \tdata_i[3] , \tdata_i[0] , \u_scaler_gray/n129 , 
        \u_scaler_gray/n128 , \u_scaler_gray/n127 , \u_scaler_gray/n126 , 
        \u_scaler_gray/n125 , \u_scaler_gray/n124 , \u_scaler_gray/n123 , 
        \u_scaler_gray/n122 , \u_scaler_gray/n121 , \u_scaler_gray/n120 , 
        \u_scaler_gray/n119 , \u_scaler_gray/n118 , \u_scaler_gray/n117 , 
        \u_scaler_gray/n116 , \u_scaler_gray/n115 , \tx_slowclk~O , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n462 , 
        \hdmi_clk1x_i~O , \hdmi_clk2x_i~O , \cmos_pclk~O , \jtag_inst1_TCK~O , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n335 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n334 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n333 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n332 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n331 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n330 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n329 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n328 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n327 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n326 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n325 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n324 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n323 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n322 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n321 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n320 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n319 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n318 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n317 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n461 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n460 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n459 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n458 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n457 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n456 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n455 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n454 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n453 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n452 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n451 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n450 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n449 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n448 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n447 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n446 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n445 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n444 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n443 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n442 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n441 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n440 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n439 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n438 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n437 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n436 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n435 , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n344 , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 , 
        n10591, n10592, n10593, n10594, n10595, n10596, n10597, 
        n10598, n10599, n10601, n10602, n10603, n10604, n10605, 
        n10606, n10607, n10608, \Axi_Clk~O , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n343 , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n342 , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n341 , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n340 , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n339 , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n338 , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n337 , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n336 , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n335 , 
        lcd_vs, \u_axi4_ctrl/n1469 , \u_axi4_ctrl/n317 , \u_axi4_ctrl/equal_38/n3 , 
        \u_axi4_ctrl/n336 , \u_axi4_ctrl/equal_47/n3 , \u_axi4_ctrl/n389 , 
        \u_axi4_ctrl/n405 , \u_axi4_ctrl/n1476 , \u_axi4_ctrl/n363 , \u_axi4_ctrl/n1544 , 
        \u_axi4_ctrl/n379 , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int , \u_axi4_ctrl/n316 , 
        ceg_net289, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] , 
        n7366, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] , 
        ceg_net296, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] , 
        \u_axi4_ctrl/n335 , \u_axi4_ctrl/n1612 , \u_axi4_ctrl/n1619 , 
        \u_axi4_ctrl/n387 , \u_axi4_ctrl/n369 , n7826, n7829, n7832, 
        n7835, n7838, n7841, n7844, n7847, n7850, n7853, n7856, 
        n7859, \u_axi4_ctrl/n381 , \u_axi4_ctrl/n1478 , \u_axi4_ctrl/n697 , 
        ceg_net401, \u_axi4_ctrl/n696 , \u_axi4_ctrl/n695 , \u_axi4_ctrl/n694 , 
        \u_axi4_ctrl/n693 , \u_axi4_ctrl/n692 , \u_axi4_ctrl/n691 , \u_axi4_ctrl/n690 , 
        \u_axi4_ctrl/n689 , \u_axi4_ctrl/n688 , \u_axi4_ctrl/n687 , \u_axi4_ctrl/n686 , 
        \u_axi4_ctrl/n685 , \u_axi4_ctrl/n684 , \u_axi4_ctrl/n683 , \u_axi4_ctrl/n682 , 
        \u_axi4_ctrl/n1499 , \u_axi4_ctrl/n1504 , \u_axi4_ctrl/n1509 , 
        \u_axi4_ctrl/n1514 , \u_axi4_ctrl/n1519 , \u_axi4_ctrl/n1524 , 
        \u_axi4_ctrl/n1529 , \u_axi4_ctrl/n1534 , \u_axi4_ctrl/n1549 , 
        \u_axi4_ctrl/n1554 , \u_axi4_ctrl/n1559 , \u_axi4_ctrl/n1564 , 
        \u_axi4_ctrl/n1569 , \u_axi4_ctrl/n1574 , \u_axi4_ctrl/n1579 , 
        \u_lcd_driver/n83 , \u_lcd_driver/equal_17/n23 , \u_lcd_driver/n35 , 
        n8110, \u_lcd_driver/n97 , \u_lcd_driver/n125 , \lcd_data[0] , 
        \u_lcd_driver/n133 , \u_lcd_driver/n34 , \u_lcd_driver/n82 , \u_lcd_driver/n81 , 
        \u_lcd_driver/n80 , \u_lcd_driver/n79 , \u_lcd_driver/n78 , \u_lcd_driver/n77 , 
        \u_lcd_driver/n76 , \u_lcd_driver/n75 , \u_lcd_driver/n74 , \u_lcd_driver/n73 , 
        \u_lcd_driver/n72 , \lcd_data[1] , \lcd_data[2] , \lcd_data[3] , 
        \lcd_data[4] , \lcd_data[5] , \lcd_data[6] , \lcd_data[7] , 
        \u_lcd_driver/n33 , \u_lcd_driver/n32 , \u_lcd_driver/n31 , \u_lcd_driver/n30 , 
        \u_lcd_driver/n29 , \u_lcd_driver/n28 , \u_lcd_driver/n27 , \u_lcd_driver/n26 , 
        \u_lcd_driver/n25 , \u_lcd_driver/n24 , \u_lcd_driver/n23 , \u_rgb2dvi/enc_0/n866 , 
        \u_rgb2dvi/enc_0/n768 , \u_rgb2dvi/enc_0/n774 , \u_rgb2dvi/enc_0/n780 , 
        \u_rgb2dvi/enc_0/n786 , \u_rgb2dvi/enc_0/n792 , \u_rgb2dvi/enc_0/n798 , 
        \u_rgb2dvi/enc_0/n804 , \u_rgb2dvi/enc_0/n810 , \u_rgb2dvi/enc_0/n816 , 
        \u_rgb2dvi/enc_1/q_out[0] , \u_rgb2dvi/enc_1/q_out[1] , \u_rgb2dvi/enc_1/q_out[2] , 
        \u_rgb2dvi/enc_1/q_out[3] , \u_rgb2dvi/enc_1/q_out[4] , \u_rgb2dvi/enc_1/q_out[5] , 
        \u_rgb2dvi/enc_1/q_out[6] , \u_rgb2dvi/enc_1/q_out[7] , \u_rgb2dvi/enc_1/q_out[9] , 
        n8411, \u_rgb2dvi/enc_2/q_out[0] , \u_rgb2dvi/enc_2/q_out[1] , 
        \u_rgb2dvi/enc_2/q_out[2] , \u_rgb2dvi/enc_2/q_out[3] , \u_rgb2dvi/enc_2/q_out[4] , 
        \u_rgb2dvi/enc_2/q_out[5] , \u_rgb2dvi/enc_2/q_out[6] , \u_rgb2dvi/enc_2/q_out[7] , 
        \u_rgb2dvi/enc_2/q_out[9] , \r_hdmi_txc_o[9] , n591, n590, n589, 
        n588, n613, n612, n611, n610, \edb_top_inst/edb_user_dr[62] , 
        \edb_top_inst/edb_user_dr[63] , \edb_top_inst/la0/n1317 , \edb_top_inst/ceg_net5 , 
        \edb_top_inst/edb_user_dr[60] , \edb_top_inst/la0/n6737 , \edb_top_inst/la0/n1318 , 
        \edb_top_inst/la0/n1319 , \edb_top_inst/edb_user_dr[0] , \edb_top_inst/la0/n1373 , 
        \edb_top_inst/edb_user_dr[42] , \edb_top_inst/la0/n1890 , \edb_top_inst/edb_user_dr[59] , 
        \edb_top_inst/la0/n1942 , \edb_top_inst/la0/data_to_addr_counter[0] , 
        \edb_top_inst/la0/addr_ct_en , \edb_top_inst/edb_user_dr[77] , \edb_top_inst/la0/op_reg_en , 
        \edb_top_inst/la0/n2166 , \edb_top_inst/ceg_net26 , \edb_top_inst/la0/data_to_word_counter[0] , 
        \edb_top_inst/la0/word_ct_en , \edb_top_inst/la0/n2443 , \edb_top_inst/ceg_net14 , 
        \edb_top_inst/la0/module_next_state[0] , \edb_top_inst/la0/n2730 , 
        \edb_top_inst/edb_user_dr[2] , \edb_top_inst/la0/n2743 , \edb_top_inst/edb_user_dr[1] , 
        \edb_top_inst/la0/n3576 , \edb_top_inst/la0/n4465 , \edb_top_inst/la0/n4480 , 
        \edb_top_inst/la0/n4678 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/edb_user_dr[64] , \edb_top_inst/la0/regsel_ld_en , 
        \edb_top_inst/edb_user_dr[43] , \edb_top_inst/edb_user_dr[61] , 
        \edb_top_inst/edb_user_dr[3] , \edb_top_inst/edb_user_dr[4] , \edb_top_inst/edb_user_dr[5] , 
        \edb_top_inst/edb_user_dr[6] , \edb_top_inst/edb_user_dr[7] , \edb_top_inst/edb_user_dr[8] , 
        \edb_top_inst/edb_user_dr[9] , \edb_top_inst/edb_user_dr[10] , \edb_top_inst/edb_user_dr[11] , 
        \edb_top_inst/edb_user_dr[12] , \edb_top_inst/edb_user_dr[13] , 
        \edb_top_inst/edb_user_dr[14] , \edb_top_inst/edb_user_dr[15] , 
        \edb_top_inst/edb_user_dr[16] , \edb_top_inst/edb_user_dr[17] , 
        \edb_top_inst/edb_user_dr[18] , \edb_top_inst/edb_user_dr[19] , 
        \edb_top_inst/edb_user_dr[20] , \edb_top_inst/edb_user_dr[21] , 
        \edb_top_inst/edb_user_dr[22] , \edb_top_inst/edb_user_dr[23] , 
        \edb_top_inst/edb_user_dr[24] , \edb_top_inst/edb_user_dr[25] , 
        \edb_top_inst/edb_user_dr[26] , \edb_top_inst/edb_user_dr[27] , 
        \edb_top_inst/edb_user_dr[28] , \edb_top_inst/edb_user_dr[29] , 
        \edb_top_inst/edb_user_dr[30] , \edb_top_inst/edb_user_dr[31] , 
        \edb_top_inst/edb_user_dr[32] , \edb_top_inst/edb_user_dr[33] , 
        \edb_top_inst/edb_user_dr[34] , \edb_top_inst/edb_user_dr[35] , 
        \edb_top_inst/edb_user_dr[36] , \edb_top_inst/edb_user_dr[37] , 
        \edb_top_inst/edb_user_dr[38] , \edb_top_inst/edb_user_dr[39] , 
        \edb_top_inst/edb_user_dr[40] , \edb_top_inst/edb_user_dr[41] , 
        \edb_top_inst/edb_user_dr[44] , \edb_top_inst/edb_user_dr[45] , 
        \edb_top_inst/edb_user_dr[46] , \edb_top_inst/edb_user_dr[47] , 
        \edb_top_inst/edb_user_dr[48] , \edb_top_inst/edb_user_dr[49] , 
        \edb_top_inst/edb_user_dr[50] , \edb_top_inst/edb_user_dr[51] , 
        \edb_top_inst/edb_user_dr[52] , \edb_top_inst/edb_user_dr[53] , 
        \edb_top_inst/edb_user_dr[54] , \edb_top_inst/edb_user_dr[55] , 
        \edb_top_inst/edb_user_dr[56] , \edb_top_inst/edb_user_dr[57] , 
        \edb_top_inst/edb_user_dr[58] , \edb_top_inst/la0/data_to_addr_counter[1] , 
        \edb_top_inst/la0/data_to_addr_counter[2] , \edb_top_inst/la0/data_to_addr_counter[3] , 
        \edb_top_inst/la0/data_to_addr_counter[4] , \edb_top_inst/la0/data_to_addr_counter[5] , 
        \edb_top_inst/la0/data_to_addr_counter[6] , \edb_top_inst/la0/data_to_addr_counter[7] , 
        \edb_top_inst/la0/data_to_addr_counter[8] , \edb_top_inst/la0/data_to_addr_counter[9] , 
        \edb_top_inst/la0/data_to_addr_counter[10] , \edb_top_inst/la0/data_to_addr_counter[11] , 
        \edb_top_inst/la0/data_to_addr_counter[12] , \edb_top_inst/la0/data_to_addr_counter[13] , 
        \edb_top_inst/la0/data_to_addr_counter[14] , \edb_top_inst/la0/data_to_addr_counter[15] , 
        \edb_top_inst/la0/data_to_addr_counter[16] , \edb_top_inst/la0/data_to_addr_counter[17] , 
        \edb_top_inst/la0/data_to_addr_counter[18] , \edb_top_inst/la0/data_to_addr_counter[19] , 
        \edb_top_inst/la0/data_to_addr_counter[20] , \edb_top_inst/la0/data_to_addr_counter[21] , 
        \edb_top_inst/la0/data_to_addr_counter[22] , \edb_top_inst/la0/data_to_addr_counter[23] , 
        \edb_top_inst/la0/data_to_addr_counter[24] , \edb_top_inst/la0/data_to_addr_counter[25] , 
        \edb_top_inst/la0/data_to_addr_counter[26] , \edb_top_inst/edb_user_dr[78] , 
        \edb_top_inst/edb_user_dr[79] , \edb_top_inst/edb_user_dr[80] , 
        \edb_top_inst/la0/n2165 , \edb_top_inst/la0/n2164 , \edb_top_inst/la0/n2163 , 
        \edb_top_inst/la0/n2162 , \edb_top_inst/la0/n2161 , \edb_top_inst/la0/data_to_word_counter[1] , 
        \edb_top_inst/la0/data_to_word_counter[2] , \edb_top_inst/la0/data_to_word_counter[3] , 
        \edb_top_inst/la0/data_to_word_counter[4] , \edb_top_inst/la0/data_to_word_counter[5] , 
        \edb_top_inst/la0/data_to_word_counter[6] , \edb_top_inst/la0/data_to_word_counter[7] , 
        \edb_top_inst/la0/data_to_word_counter[8] , \edb_top_inst/la0/data_to_word_counter[9] , 
        \edb_top_inst/la0/data_to_word_counter[10] , \edb_top_inst/la0/data_to_word_counter[11] , 
        \edb_top_inst/la0/data_to_word_counter[12] , \edb_top_inst/la0/data_to_word_counter[13] , 
        \edb_top_inst/la0/data_to_word_counter[14] , \edb_top_inst/la0/data_to_word_counter[15] , 
        \edb_top_inst/la0/n2442 , \edb_top_inst/la0/n2441 , \edb_top_inst/la0/n2440 , 
        \edb_top_inst/la0/n2439 , \edb_top_inst/la0/n2438 , \edb_top_inst/la0/n2437 , 
        \edb_top_inst/la0/n2436 , \edb_top_inst/la0/n2435 , \edb_top_inst/la0/n2434 , 
        \edb_top_inst/la0/n2433 , \edb_top_inst/la0/n2432 , \edb_top_inst/la0/n2431 , 
        \edb_top_inst/la0/n2430 , \edb_top_inst/la0/n2429 , \edb_top_inst/la0/n2428 , 
        \edb_top_inst/la0/n2427 , \edb_top_inst/la0/n2426 , \edb_top_inst/la0/n2425 , 
        \edb_top_inst/la0/n2424 , \edb_top_inst/la0/n2423 , \edb_top_inst/la0/n2422 , 
        \edb_top_inst/la0/n2421 , \edb_top_inst/la0/n2420 , \edb_top_inst/la0/n2419 , 
        \edb_top_inst/la0/n2418 , \edb_top_inst/la0/n2417 , \edb_top_inst/la0/n2416 , 
        \edb_top_inst/la0/n2415 , \edb_top_inst/la0/n2414 , \edb_top_inst/la0/n2413 , 
        \edb_top_inst/la0/n2412 , \edb_top_inst/la0/n2411 , \edb_top_inst/la0/n2410 , 
        \edb_top_inst/la0/n2409 , \edb_top_inst/la0/n2408 , \edb_top_inst/la0/n2407 , 
        \edb_top_inst/la0/n2406 , \edb_top_inst/la0/n2405 , \edb_top_inst/la0/n2404 , 
        \edb_top_inst/la0/n2403 , \edb_top_inst/la0/n2402 , \edb_top_inst/la0/n2401 , 
        \edb_top_inst/la0/n2400 , \edb_top_inst/la0/n2399 , \edb_top_inst/la0/n2398 , 
        \edb_top_inst/la0/n2397 , \edb_top_inst/la0/n2396 , \edb_top_inst/la0/n2395 , 
        \edb_top_inst/la0/n2394 , \edb_top_inst/la0/n2393 , \edb_top_inst/la0/n2392 , 
        \edb_top_inst/la0/n2391 , \edb_top_inst/la0/n2390 , \edb_top_inst/la0/n2389 , 
        \edb_top_inst/la0/n2388 , \edb_top_inst/la0/n2387 , \edb_top_inst/la0/n2386 , 
        \edb_top_inst/la0/n2385 , \edb_top_inst/la0/n2384 , \edb_top_inst/la0/n2383 , 
        \edb_top_inst/la0/n2382 , \edb_top_inst/la0/n2381 , \edb_top_inst/la0/n2380 , 
        \edb_top_inst/la0/module_next_state[1] , \edb_top_inst/la0/module_next_state[2] , 
        \edb_top_inst/la0/module_next_state[3] , \edb_top_inst/la0/axi_crc_i/n150 , 
        \edb_top_inst/ceg_net221 , \edb_top_inst/la0/axi_crc_i/n149 , \edb_top_inst/la0/axi_crc_i/n148 , 
        \edb_top_inst/la0/axi_crc_i/n147 , \edb_top_inst/la0/axi_crc_i/n146 , 
        \edb_top_inst/la0/axi_crc_i/n145 , \edb_top_inst/la0/axi_crc_i/n144 , 
        \edb_top_inst/la0/axi_crc_i/n143 , \edb_top_inst/la0/axi_crc_i/n142 , 
        \edb_top_inst/la0/axi_crc_i/n141 , \edb_top_inst/la0/axi_crc_i/n140 , 
        \edb_top_inst/la0/axi_crc_i/n139 , \edb_top_inst/la0/axi_crc_i/n138 , 
        \edb_top_inst/la0/axi_crc_i/n137 , \edb_top_inst/la0/axi_crc_i/n136 , 
        \edb_top_inst/la0/axi_crc_i/n135 , \edb_top_inst/la0/axi_crc_i/n134 , 
        \edb_top_inst/la0/axi_crc_i/n133 , \edb_top_inst/la0/axi_crc_i/n132 , 
        \edb_top_inst/la0/axi_crc_i/n131 , \edb_top_inst/la0/axi_crc_i/n130 , 
        \edb_top_inst/la0/axi_crc_i/n129 , \edb_top_inst/la0/axi_crc_i/n128 , 
        \edb_top_inst/la0/axi_crc_i/n127 , \edb_top_inst/la0/axi_crc_i/n126 , 
        \edb_top_inst/la0/axi_crc_i/n125 , \edb_top_inst/la0/axi_crc_i/n124 , 
        \edb_top_inst/la0/axi_crc_i/n123 , \edb_top_inst/la0/axi_crc_i/n122 , 
        \edb_top_inst/la0/axi_crc_i/n121 , \edb_top_inst/la0/axi_crc_i/n120 , 
        \edb_top_inst/la0/axi_crc_i/n119 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n19 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n16 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n17 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n19 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n41 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n50 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n39 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n38 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n37 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n36 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n35 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n34 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n33 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n21 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n20 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n19 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n15 , \edb_top_inst/la0/trigger_tu/n35 , 
        \edb_top_inst/la0/la_biu_inst/next_state[0] , \edb_top_inst/la0/la_biu_inst/run_trig_p1 , 
        \edb_top_inst/la0/la_biu_inst/n350 , \edb_top_inst/la0/la_biu_inst/n1251 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[0] , \edb_top_inst/la0/la_biu_inst/next_fsm_state[0] , 
        \edb_top_inst/ceg_net351 , \edb_top_inst/la0/la_biu_inst/n1236 , 
        \edb_top_inst/la0/n7224 , \edb_top_inst/la0/la_biu_inst/next_state[2] , 
        \edb_top_inst/la0/la_biu_inst/next_state[1] , \edb_top_inst/ceg_net348 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[1] , \edb_top_inst/la0/la_biu_inst/fifo_dout[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[3] , \edb_top_inst/la0/la_biu_inst/fifo_dout[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[5] , \edb_top_inst/la0/la_biu_inst/fifo_dout[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[7] , \edb_top_inst/la0/la_biu_inst/fifo_dout[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[9] , \edb_top_inst/la0/la_biu_inst/fifo_dout[10] , 
        \edb_top_inst/la0/la_biu_inst/next_fsm_state[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data , 
        \edb_top_inst/la0/la_biu_inst/fifo_rstn , \edb_top_inst/la0/la_biu_inst/n1993 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 , \edb_top_inst/la0/la_biu_inst/fifo_push , 
        \edb_top_inst/ceg_net355 , \edb_top_inst/n297 , \edb_top_inst/n765 , 
        \edb_top_inst/n763 , \edb_top_inst/n761 , \edb_top_inst/n759 , 
        \edb_top_inst/n757 , \edb_top_inst/n755 , \edb_top_inst/n753 , 
        \edb_top_inst/n751 , \edb_top_inst/n749 , \edb_top_inst/n748 , 
        \edb_top_inst/n426 , \edb_top_inst/n746 , \edb_top_inst/n744 , 
        \edb_top_inst/n742 , \edb_top_inst/n740 , \edb_top_inst/n738 , 
        \edb_top_inst/n736 , \edb_top_inst/n734 , \edb_top_inst/n732 , 
        \edb_top_inst/n730 , \edb_top_inst/n727 , \edb_top_inst/n428 , 
        \edb_top_inst/n695 , \edb_top_inst/n693 , \edb_top_inst/n691 , 
        \edb_top_inst/n689 , \edb_top_inst/n687 , \edb_top_inst/n685 , 
        \edb_top_inst/n683 , \edb_top_inst/n681 , \edb_top_inst/n679 , 
        \edb_top_inst/n677 , \edb_top_inst/n434 , \edb_top_inst/n630 , 
        \edb_top_inst/n628 , \edb_top_inst/n626 , \edb_top_inst/n624 , 
        \edb_top_inst/n622 , \edb_top_inst/n620 , \edb_top_inst/n618 , 
        \edb_top_inst/n616 , \edb_top_inst/n614 , \edb_top_inst/n612 , 
        \edb_top_inst/n590 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] , 
        \edb_top_inst/n432 , \edb_top_inst/n651 , \edb_top_inst/n649 , 
        \edb_top_inst/n647 , \edb_top_inst/n645 , \edb_top_inst/n643 , 
        \edb_top_inst/n641 , \edb_top_inst/n639 , \edb_top_inst/n637 , 
        \edb_top_inst/n635 , \edb_top_inst/n633 , \edb_top_inst/n632 , 
        \edb_top_inst/edb_user_dr[65] , \edb_top_inst/edb_user_dr[66] , 
        \edb_top_inst/edb_user_dr[67] , \edb_top_inst/edb_user_dr[68] , 
        \edb_top_inst/edb_user_dr[69] , \edb_top_inst/edb_user_dr[70] , 
        \edb_top_inst/edb_user_dr[71] , \edb_top_inst/edb_user_dr[72] , 
        \edb_top_inst/edb_user_dr[73] , \edb_top_inst/edb_user_dr[74] , 
        \edb_top_inst/edb_user_dr[75] , \edb_top_inst/edb_user_dr[76] , 
        \edb_top_inst/debug_hub_inst/n266 , \edb_top_inst/debug_hub_inst/n95 , 
        \edb_top_inst/edb_user_dr[81] , \edb_top_inst/n613 , \edb_top_inst/n615 , 
        \edb_top_inst/n617 , \edb_top_inst/n619 , \edb_top_inst/n621 , 
        \edb_top_inst/n623 , \edb_top_inst/n625 , \edb_top_inst/n627 , 
        \edb_top_inst/n629 , \edb_top_inst/n631 , \edb_top_inst/n634 , 
        \edb_top_inst/n636 , \edb_top_inst/n638 , \edb_top_inst/n640 , 
        \edb_top_inst/n642 , \edb_top_inst/n644 , \edb_top_inst/n646 , 
        \edb_top_inst/n648 , \edb_top_inst/n650 , \edb_top_inst/n652 , 
        \edb_top_inst/n680 , \edb_top_inst/n682 , \edb_top_inst/n684 , 
        \edb_top_inst/n686 , \edb_top_inst/n688 , \edb_top_inst/n690 , 
        \edb_top_inst/n692 , \edb_top_inst/n694 , \edb_top_inst/n696 , 
        \edb_top_inst/n731 , \edb_top_inst/n733 , \edb_top_inst/n735 , 
        \edb_top_inst/n737 , \edb_top_inst/n739 , \edb_top_inst/n741 , 
        \edb_top_inst/n743 , \edb_top_inst/n745 , \edb_top_inst/n747 , 
        \edb_top_inst/n750 , \edb_top_inst/n752 , \edb_top_inst/n754 , 
        \edb_top_inst/n756 , \edb_top_inst/n758 , \edb_top_inst/n760 , 
        \edb_top_inst/n762 , \edb_top_inst/n764 , \edb_top_inst/n766 , 
        \edb_top_inst/n769 , \edb_top_inst/n771 , \edb_top_inst/n773 , 
        \edb_top_inst/n786 , \edb_top_inst/n788 , \edb_top_inst/n790 , 
        \edb_top_inst/n792 , \edb_top_inst/n794 , \edb_top_inst/n796 , 
        \edb_top_inst/n798 , \edb_top_inst/n800 , \edb_top_inst/n802 , 
        \edb_top_inst/n804 , \edb_top_inst/n806 , \edb_top_inst/n808 , 
        \edb_top_inst/n810 , \edb_top_inst/n812 , \edb_top_inst/n814 , 
        \edb_top_inst/n816 , \edb_top_inst/n818 , \edb_top_inst/n820 , 
        \edb_top_inst/n822 , \edb_top_inst/n824 , \edb_top_inst/n826 , 
        \edb_top_inst/n828 , \edb_top_inst/n830 , \edb_top_inst/n832 , 
        \edb_top_inst/n834 , \edb_top_inst/n847 , \edb_top_inst/n849 , 
        \edb_top_inst/n851 , \edb_top_inst/n853 , \edb_top_inst/n855 , 
        \edb_top_inst/n857 , \edb_top_inst/n862 , \edb_top_inst/n864 , 
        \edb_top_inst/n866 , \edb_top_inst/n868 , \edb_top_inst/n1730 , 
        \edb_top_inst/n34 , \edb_top_inst/n833 , \edb_top_inst/n831 , 
        \edb_top_inst/n829 , \edb_top_inst/n827 , \edb_top_inst/n825 , 
        \edb_top_inst/n823 , \edb_top_inst/n821 , \edb_top_inst/n819 , 
        \edb_top_inst/n817 , \edb_top_inst/n815 , \edb_top_inst/n813 , 
        \edb_top_inst/n811 , \edb_top_inst/n809 , \edb_top_inst/n807 , 
        \edb_top_inst/n805 , \edb_top_inst/n803 , \edb_top_inst/n867 , 
        \edb_top_inst/n801 , \edb_top_inst/n865 , \edb_top_inst/n799 , 
        \edb_top_inst/n863 , \edb_top_inst/n797 , \edb_top_inst/n861 , 
        \edb_top_inst/n795 , \edb_top_inst/n856 , \edb_top_inst/n793 , 
        \edb_top_inst/n854 , \edb_top_inst/n791 , \edb_top_inst/n852 , 
        \edb_top_inst/n789 , \edb_top_inst/n850 , \edb_top_inst/n787 , 
        \edb_top_inst/n848 , \edb_top_inst/n785 , \edb_top_inst/n846 , 
        \edb_top_inst/n783 , \edb_top_inst/n844 , \edb_top_inst/n36 , 
        \edb_top_inst/n772 , \edb_top_inst/n770 , \edb_top_inst/n768 , 
        \edb_top_inst/n767 , \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q_pinv , 
        \u_lcd_driver/vcnt[7]~FF_frt_39_q_pinv , \u_lcd_driver/vcnt[2]~FF_frt_40_q_pinv , 
        \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q_pinv , \u_lcd_driver/hcnt[8]~FF_frt_41_q , 
        \u_lcd_driver/vcnt[2]~FF_frt_40_q , \u_lcd_driver/vcnt[7]~FF_frt_39_q , 
        \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38_q , \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q , 
        \u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36_q , \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35_q , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32_q , 
        \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q , \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27_q , 
        \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26_q , \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q , 
        \u_lcd_driver/r_lcd_rgb[0]~FF_frt_24_q , \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_q , 
        \u_lcd_driver/r_lcd_rgb[0]~FF_frt_11_q , \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_q , 
        \u_lcd_driver/r_lcd_dv~FF_frt_7_q , \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3_q , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2_q , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1_q , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_q , 
        n10069, n10070, n10071, n10072, n10073, n10074, n10075, 
        n10076, n10077, n10078, n10079, n10080, n10081, n10082, 
        n10083, n10084, n10085, n10086, n10087, n10088, n10089, 
        n10090, n10091, n10092, n10093, n10094, n10095, n10096, 
        n10097, n10098, n10099, n10100, n10101, n10102, n10103, 
        n10104, n10105, n10106, n10107, n10108, n10109, n10110, 
        n10111, n10112, n10113, n10114, n10115, n10116, n10117, 
        n10118, n10119, n10120, n10121, n10122, n10123, n10124, 
        n10125, n10126, n10127, n10128, n10129, n10130, n10131, 
        n10132, n10133, n10134, n10135, n10136, n10137, n10138, 
        n10139, n10140, n10141, n10142, n10143, n10144, n10145, 
        n10146, n10147, n10148, n10149, n10150, n10151, n10152, 
        n10153, n10154, n10155, n10156, n10157, n10158, n10159, 
        n10160, n10161, n10162, n10163, n10164, n10165, n10166, 
        n10167, n10168, n10169, n10170, n10171, n10172, n10173, 
        n10174, n10175, n10176, n10177, n10178, n10179, n10180, 
        n10181, n10182, n10183, n10184, n10185, n10186, n10187, 
        n10188, n10189, n10190, n10191, n10192, n10193, n10194, 
        n10195, n10196, n10197, n10198, n10199, n10200, n10201, 
        n10202, n10203, n10204, n10205, n10206, n10207, n10208, 
        n10209, n10210, n10211, n10212, n10213, n10214, n10215, 
        n10216, n10217, n10218, n10219, n10220, n10221, n10222, 
        n10223, n10224, n10225, n10226, n10227, n10228, n10229, 
        n10230, n10231, n10232, n10233, n10234, n10235, n10236, 
        n10237, n10238, n10239, n10240, n10241, n10242, n10243, 
        n10244, n10245, n10246, n10247, n10248, n10249, n10250, 
        n10251, n10252, n10253, n10254, n10255, n10256, n10257, 
        n10258, n10259, n10260, n10261, n10262, n10263, n10264, 
        n10265, n10266, n10267, n10268, n10269, n10270, n10271, 
        n10272, n10273, n10274, n10275, n10276, n10277, n10278, 
        n10279, n10280, n10281, n10282, n10283, n10284, n10285, 
        n10286, n10287, n10288, n10289, n10290, n10291, n10292, 
        n10293, n10294, n10295, n10296, n10297, n10298, n10299, 
        n10300, n10301, n10302, n10303, n10304, n10305, n10306, 
        n10307, n10308, n10309, n10310, n10311, n10312, n10313, 
        n10314, n10315, n10316, n10317, n10318, n10319, n10320, 
        n10321, n10322, n10323, n10324, n10325, n10326, n10327, 
        n10330, n10347, n10348, n10349, n10350, n10351, n10352, 
        n10353, n10354, n10355, n10356, n10357, n10358, n10359, 
        n10360, n10361, n10362, n10363, n10364, n10365, n10366, 
        n10367, n10368, n10369, n10370, n10371, n10372, n10373, 
        n10374, n10375, n10376, n10377, n10378, n10379, n10380, 
        n10381, n10382, n10383, n10384, n10385, n10386, n10387, 
        n10388, n10389, n10390, n10391, n10392, n10393, n10394, 
        n10395, n10396, n10397, n10398, n10399, n10400, n10401, 
        n10402, n10403, n10404, n10405, n10406, n10407, n10408, 
        n10409, n10410, n10411, n10412, n10413, n10414, n10415, 
        n10416, n10417, n10418, n10419, n10420, n10421, n10422, 
        n10423, n10424, n10425, n10426, n10427, n10428, n10429, 
        n10430, n10431, n10432, n10433, n10434, n10435, n10436, 
        n10437, n10438, n10439, n10440, n10441, n10442, n10443, 
        n10444, n10445, n10446, n10447, n10448, n10449, n10450, 
        n10451, n10452, n10453, n10454, n10455, n10456, n10457, 
        n10458, n10459, n10460, n10461, n10462, n10463, n10464, 
        n10465, n10466, n10467, n10468, n10469, n10470, n10471, 
        n10472, n10473, n10474, n10475, n10476, n10477, n10478, 
        n10479, n10480, n10481, n10482, n10483, n10484, n10485, 
        n10486, n10487, n10488, n10489, n10490, n10491, n10492, 
        n10493, n10494, n10495, n10496, n10497, n10498, n10499, 
        n10500, n10501, n10502, n10503, n10504, n10505, n10506, 
        n10507, n10508, n10509, n10510, n10511, n10512, n10513, 
        n10514, n10515, n10516, n10517, n10518, n10519, n10520, 
        n10521, n10524, n10525, n10526, n10527, n10528, n10529, 
        n10530, n10531, n10532, n10533, n10534, n10535, n10536, 
        n10537, n10538, n10539, n10540, n10541, n10542, n10543, 
        n10544, n10545, n10546, n10547, n10548, n10549, n10550, 
        n10551, n10552, n10553, n10554, n10555, n10556, n10557, 
        n10558, n10559, n10560, n10561, n10562, n10563, n10564, 
        n10565, n10566, n10567, n10568, n10569, n10570, n10571, 
        n10572, n10573, n10574, n10575, n10576, n10577, n10578, 
        n10579, n10580, n10581, n10582, n10583, n10584, n10585, 
        n10586, n10587, n10588, n10589, n10590;
    
    assign DdrCtrl_AID_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[31] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[30] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[29] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[28] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[27] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[26] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[9] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[8] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[5] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[4] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[3] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[2] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[1] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[2] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ABURST_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ABURST_0[0] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALOCK_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALOCK_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[15] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[14] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[13] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[12] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[11] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[10] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[9] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[8] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[7] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[6] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[5] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[4] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[3] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[2] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[1] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[0] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign cmos_ctl0 = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign cmos_ctl2 = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign cmos_ctl3 = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[4] = hdmi_txc_o[2] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[3] = hdmi_txc_o[2] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[1] = hdmi_txc_o[2] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[0] = hdmi_txc_o[2] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lcd_pwm = 1'b1 /* verific EFX_ATTRIBUTE_CELL_NAME=VCC */ ;
    assign lvds_tx0_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_LUT4 \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_rtinv  (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q_pinv ), 
            .O(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_rtinv .LUTMASK = 16'h5555;
    EFX_FF \ResetShiftReg[0]~FF  (.D(\reduce_nand_9/n7 ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\ResetShiftReg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(128)
    defparam \ResetShiftReg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .CE_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .D_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_SYNC = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_VALUE = 1'b0;
    defparam \ResetShiftReg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[0]~FF  (.D(DdrInitDone), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(161)
    defparam \Axi0ResetReg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_rst_n~FF  (.D(\Axi0ResetReg[2] ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(r_hdmi_rst_n)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(456)
    defparam \r_hdmi_rst_n~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .SR_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_rst_n~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_rst_n~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rc_hdmi_tx~FF  (.D(rc_hdmi_tx), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(rc_hdmi_tx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \rc_hdmi_tx~FF .CLK_POLARITY = 1'b1;
    defparam \rc_hdmi_tx~FF .CE_POLARITY = 1'b1;
    defparam \rc_hdmi_tx~FF .SR_POLARITY = 1'b1;
    defparam \rc_hdmi_tx~FF .D_POLARITY = 1'b0;
    defparam \rc_hdmi_tx~FF .SR_SYNC = 1'b1;
    defparam \rc_hdmi_tx~FF .SR_VALUE = 1'b0;
    defparam \rc_hdmi_tx~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[0]~FF  (.D(n592_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx0_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[0]~FF  (.D(n603_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx1_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[0]~FF  (.D(n614_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx2_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[0]~FF  (.D(n4990), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ResetShiftReg[1]~FF  (.D(\ResetShiftReg[0] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\ResetShiftReg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(128)
    defparam \ResetShiftReg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .CE_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .D_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_SYNC = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_VALUE = 1'b0;
    defparam \ResetShiftReg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_CFG_RST_N~FF  (.D(\ResetShiftReg[1] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(DdrCtrl_CFG_RST_N)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(128)
    defparam \DdrCtrl_CFG_RST_N~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[1]~FF  (.D(\Axi0ResetReg[0] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(161)
    defparam \Axi0ResetReg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[2]~FF  (.D(\Axi0ResetReg[1] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(161)
    defparam \Axi0ResetReg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrInitDone~FF  (.D(1'b1), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(DdrInitDone)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \DdrInitDone~FF .CLK_POLARITY = 1'b1;
    defparam \DdrInitDone~FF .CE_POLARITY = 1'b0;
    defparam \DdrInitDone~FF .SR_POLARITY = 1'b0;
    defparam \DdrInitDone~FF .D_POLARITY = 1'b1;
    defparam \DdrInitDone~FF .SR_SYNC = 1'b0;
    defparam \DdrInitDone~FF .SR_VALUE = 1'b0;
    defparam \DdrInitDone~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_CFG_SEQ_START~FF  (.D(1'b1), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/equal_21/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(DdrCtrl_CFG_SEQ_START)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(186)
    defparam \DdrCtrl_CFG_SEQ_START~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_SEQ_START~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n92 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(186)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(150)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF  (.D(n186), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n91 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(186)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(150)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF  (.D(n3433), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF  (.D(n3431), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF  (.D(n3429), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF  (.D(n3427), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF  (.D(n3425), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF  (.D(n3423), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF  (.D(n3421), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF  (.D(n3419), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF  (.D(n3417), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF  (.D(n3415), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF  (.D(n3413), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF  (.D(n3411), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF  (.D(n3409), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF  (.D(n3407), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF  (.D(n3405), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF  (.D(n3403), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF  (.D(n3401), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF  (.D(n3399), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF  (.D(n3398), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n137 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(167)
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n138 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n139 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n140 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n205 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[0]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[0]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[0]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[0]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n500 ), 
           .CE(ceg_net552), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n509 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n567 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n570 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n573 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n576 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n579 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n581 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF  (.D(n205), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cmos_sdat_OUT~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n495 ), .CE(ceg_net632), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(cmos_sdat_OUT)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \cmos_sdat_OUT~FF .CLK_POLARITY = 1'b1;
    defparam \cmos_sdat_OUT~FF .CE_POLARITY = 1'b1;
    defparam \cmos_sdat_OUT~FF .SR_POLARITY = 1'b0;
    defparam \cmos_sdat_OUT~FF .D_POLARITY = 1'b1;
    defparam \cmos_sdat_OUT~FF .SR_SYNC = 1'b0;
    defparam \cmos_sdat_OUT~FF .SR_VALUE = 1'b1;
    defparam \cmos_sdat_OUT~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n136 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n135 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n134 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n133 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n132 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n131 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n130 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n129 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n128 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n127 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n126 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n125 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n124 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n123 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n122 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(167)
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(167)
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(167)
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(167)
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[1]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n204 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[1]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[1]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[1]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[1]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[2]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n203 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[2]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[2]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[2]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[2]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[3]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n202 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[3]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[3]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[3]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[3]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[4]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n201 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[4]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[4]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[4]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[4]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[5]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n200 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[5]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[5]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[5]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[5]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[6]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n199 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[6]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[6]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[6]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[6]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[7]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n198 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[7]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[7]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[7]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[7]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n499 ), 
           .CE(ceg_net552), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n498 ), 
           .CE(ceg_net552), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n497 ), 
           .CE(ceg_net552), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n508 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n507 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n506 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n505 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n504 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n503 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n502 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF  (.D(n3392), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF  (.D(n3390), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF  (.D(n3388), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF  (.D(n3386), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF  (.D(n3384), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF  (.D(n3382), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF  (.D(n3380), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF  (.D(n3378), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF  (.D(n3368), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF  (.D(n3366), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF  (.D(n3364), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF  (.D(n3362), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF  (.D(n3360), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF  (.D(n3358), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF  (.D(n3356), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF  (.D(n3354), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF  (.D(n3352), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF  (.D(n3351), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF  (.D(cmos_href), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_href_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF  (.D(cmos_data[0]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n127 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n160 ), 
           .CE(ceg_net154), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(128)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF  (.D(1'b1), .CE(\u_CMOS_Capture_RAW_Gray/n171 ), 
           .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/frame_sync_flag )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(141)
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF  (.D(cmos_vsync), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_href_r[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_href_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF  (.D(cmos_data[1]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF  (.D(cmos_data[2]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF  (.D(cmos_data[3]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF  (.D(cmos_data[4]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF  (.D(cmos_data[5]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF  (.D(cmos_data[6]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF  (.D(cmos_data[7]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n126 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n125 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n124 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n123 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n122 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n121 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n120 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n119 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n118 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n117 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n116 ), 
           .CE(ceg_net126), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n159 ), 
           .CE(ceg_net154), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(128)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[0]~FF  (.D(\u_sensor_frame_count/n141 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[0]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[1] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[0]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[0]~FF .CE_POLARITY = 1'b0;
    defparam \LED[0]~FF .SR_POLARITY = 1'b0;
    defparam \LED[0]~FF .D_POLARITY = 1'b1;
    defparam \LED[0]~FF .SR_SYNC = 1'b0;
    defparam \LED[0]~FF .SR_VALUE = 1'b0;
    defparam \LED[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_vsync_r[0]~FF  (.D(cmos_vsync), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/cmos_vsync_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(53)
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[0]~FF  (.D(\u_sensor_frame_count/n75 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[1]~FF  (.D(\u_sensor_frame_count/n74 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[2]~FF  (.D(\u_sensor_frame_count/n73 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[3]~FF  (.D(\u_sensor_frame_count/n72 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[4]~FF  (.D(\u_sensor_frame_count/n71 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[5]~FF  (.D(\u_sensor_frame_count/n70 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[6]~FF  (.D(\u_sensor_frame_count/n69 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[7]~FF  (.D(\u_sensor_frame_count/n68 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[8]~FF  (.D(\u_sensor_frame_count/n67 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[9]~FF  (.D(\u_sensor_frame_count/n66 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[10]~FF  (.D(\u_sensor_frame_count/n65 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[11]~FF  (.D(\u_sensor_frame_count/n64 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[12]~FF  (.D(\u_sensor_frame_count/n63 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[13]~FF  (.D(\u_sensor_frame_count/n62 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[14]~FF  (.D(\u_sensor_frame_count/n61 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[15]~FF  (.D(\u_sensor_frame_count/n60 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[16]~FF  (.D(\u_sensor_frame_count/n59 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[17]~FF  (.D(\u_sensor_frame_count/n58 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[18]~FF  (.D(\u_sensor_frame_count/n57 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[19]~FF  (.D(\u_sensor_frame_count/n56 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[20]~FF  (.D(\u_sensor_frame_count/n55 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[21]~FF  (.D(\u_sensor_frame_count/n54 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[22]~FF  (.D(\u_sensor_frame_count/n53 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[23]~FF  (.D(\u_sensor_frame_count/n52 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[24]~FF  (.D(\u_sensor_frame_count/n51 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[25]~FF  (.D(\u_sensor_frame_count/n50 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[26]~FF  (.D(\u_sensor_frame_count/n49 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[27]~FF  (.D(\u_sensor_frame_count/n48 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[1]~FF  (.D(\u_sensor_frame_count/n140 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[2]~FF  (.D(\u_sensor_frame_count/n139 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[3]~FF  (.D(\u_sensor_frame_count/n138 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[4]~FF  (.D(\u_sensor_frame_count/n137 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[5]~FF  (.D(\u_sensor_frame_count/n136 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[6]~FF  (.D(\u_sensor_frame_count/n135 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[7]~FF  (.D(\u_sensor_frame_count/n134 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[8]~FF  (.D(\u_sensor_frame_count/n133 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[1]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[2] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[1]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[1]~FF .CE_POLARITY = 1'b0;
    defparam \LED[1]~FF .SR_POLARITY = 1'b0;
    defparam \LED[1]~FF .D_POLARITY = 1'b1;
    defparam \LED[1]~FF .SR_SYNC = 1'b0;
    defparam \LED[1]~FF .SR_VALUE = 1'b0;
    defparam \LED[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[2]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[3] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[2]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[2]~FF .CE_POLARITY = 1'b0;
    defparam \LED[2]~FF .SR_POLARITY = 1'b0;
    defparam \LED[2]~FF .D_POLARITY = 1'b1;
    defparam \LED[2]~FF .SR_SYNC = 1'b0;
    defparam \LED[2]~FF .SR_VALUE = 1'b0;
    defparam \LED[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[3]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[4] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[3]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[3]~FF .CE_POLARITY = 1'b0;
    defparam \LED[3]~FF .SR_POLARITY = 1'b0;
    defparam \LED[3]~FF .D_POLARITY = 1'b1;
    defparam \LED[3]~FF .SR_SYNC = 1'b0;
    defparam \LED[3]~FF .SR_VALUE = 1'b0;
    defparam \LED[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[4]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[5] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[4]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[4]~FF .CE_POLARITY = 1'b0;
    defparam \LED[4]~FF .SR_POLARITY = 1'b0;
    defparam \LED[4]~FF .D_POLARITY = 1'b1;
    defparam \LED[4]~FF .SR_SYNC = 1'b0;
    defparam \LED[4]~FF .SR_VALUE = 1'b0;
    defparam \LED[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[5]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[6] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[5]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[5]~FF .CE_POLARITY = 1'b0;
    defparam \LED[5]~FF .SR_POLARITY = 1'b0;
    defparam \LED[5]~FF .D_POLARITY = 1'b1;
    defparam \LED[5]~FF .SR_SYNC = 1'b0;
    defparam \LED[5]~FF .SR_VALUE = 1'b0;
    defparam \LED[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[6]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[7] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[6]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[6]~FF .CE_POLARITY = 1'b0;
    defparam \LED[6]~FF .SR_POLARITY = 1'b0;
    defparam \LED[6]~FF .D_POLARITY = 1'b1;
    defparam \LED[6]~FF .SR_SYNC = 1'b0;
    defparam \LED[6]~FF .SR_VALUE = 1'b0;
    defparam \LED[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[7]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[8] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[7]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[7]~FF .CE_POLARITY = 1'b0;
    defparam \LED[7]~FF .SR_POLARITY = 1'b0;
    defparam \LED[7]~FF .D_POLARITY = 1'b1;
    defparam \LED[7]~FF .SR_SYNC = 1'b0;
    defparam \LED[7]~FF .SR_VALUE = 1'b0;
    defparam \LED[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_vsync_r[1]~FF  (.D(\u_sensor_frame_count/cmos_vsync_r[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/cmos_vsync_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(53)
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(499)
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF  (.D(1'b0), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(499)
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF  (.D(1'b0), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(492)
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(721)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/waddr[0] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), .CLK(\cmos_pclk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/waddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \empty~FF  (.D(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CE(ceg_net219), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(empty)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1090)
    defparam \empty~FF .CLK_POLARITY = 1'b1;
    defparam \empty~FF .CE_POLARITY = 1'b0;
    defparam \empty~FF .SR_POLARITY = 1'b1;
    defparam \empty~FF .D_POLARITY = 1'b0;
    defparam \empty~FF .SR_SYNC = 1'b0;
    defparam \empty~FF .SR_VALUE = 1'b1;
    defparam \empty~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/raddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF  (.D(n694), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF  (.D(n713), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF  (.D(n2821), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF  (.D(n2819), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF  (.D(n2817), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF  (.D(n2815), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF  (.D(n2813), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF  (.D(n2811), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF  (.D(n2809), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF  (.D(n2807), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF  (.D(n2805), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF  (.D(n2803), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF  (.D(n2802), 
           .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), .CLK(\cmos_pclk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF  (.D(n719), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF  (.D(n2786), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF  (.D(n2784), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF  (.D(n2782), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF  (.D(n2780), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF  (.D(n2778), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF  (.D(n2776), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF  (.D(n2774), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF  (.D(n2772), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF  (.D(n2770), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF  (.D(n2768), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF  (.D(n2766), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF  (.D(n2765), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[1] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[2] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[3] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[4] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[5] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[6] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[7] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[8] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[9] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[10] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[11] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[13] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[12] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4  (.D(n10279), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3  (.D(n10424), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true", INIT_VALUE=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3 .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3 .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3 .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3 .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3 .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3 .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2  (.D(n10423), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true", INIT_VALUE=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1  (.D(n7829), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true", INIT_VALUE=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1 .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1 .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1 .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1 .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1 .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1 .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(492)
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[0]~FF  (.D(\u_scaler_gray/vs_cnt[0] ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tvsync_o~FF  (.D(\u_scaler_gray/n150 ), .CE(ceg_net229), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(tvsync_o)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(123)
    defparam \tvsync_o~FF .CLK_POLARITY = 1'b1;
    defparam \tvsync_o~FF .CE_POLARITY = 1'b0;
    defparam \tvsync_o~FF .SR_POLARITY = 1'b0;
    defparam \tvsync_o~FF .D_POLARITY = 1'b0;
    defparam \tvsync_o~FF .SR_SYNC = 1'b0;
    defparam \tvsync_o~FF .SR_VALUE = 1'b0;
    defparam \tvsync_o~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/tvalid_o_r~FF  (.D(tvalid_o), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\u_scaler_gray/tvalid_o_r )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(97)
    defparam \u_scaler_gray/tvalid_o_r~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid_o_r~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid_o_r~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid_o_r~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid_o_r~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/tvalid_o_r~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/tvalid_o_r~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] ), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/w_addra[0] ), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n432 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(176)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n2157 ), 
           .CE(ceg_net526), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(176)
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[0]~FF  (.D(\u_scaler_gray/destx[0] ), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[0]~FF  (.D(\u_scaler_gray/desty[0] ), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/desty[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n903 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n903 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0] ), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF  (.D(n916), .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF  (.D(n2553), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF  (.D(n2551), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF  (.D(n2549), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF  (.D(n2547), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF  (.D(n2545), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF  (.D(n2533), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF  (.D(n2528), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF  (.D(n2505), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF  (.D(n2503), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF  (.D(n2501), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF  (.D(n2499), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF  (.D(n2497), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF  (.D(n2495), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF  (.D(n2494), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF  (.D(n923), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF  (.D(n2492), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF  (.D(n2490), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF  (.D(n2488), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF  (.D(n2407), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF  (.D(n2405), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF  (.D(n2403), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF  (.D(n2401), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF  (.D(n2399), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF  (.D(n2397), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF  (.D(n2387), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF  (.D(n2385), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF  (.D(n2383), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF  (.D(n2381), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF  (.D(n2380), .CE(n197), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n431 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(176)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n430 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(176)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n2080 ), 
           .CE(ceg_net526), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(176)
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[1]~FF  (.D(n930), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[2]~FF  (.D(n2378), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[3]~FF  (.D(n2376), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[4]~FF  (.D(n2357), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[5]~FF  (.D(n2353), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[6]~FF  (.D(n2348), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[7]~FF  (.D(n2346), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[8]~FF  (.D(n2220), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[9]~FF  (.D(n2218), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[9]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[10]~FF  (.D(n2216), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[10]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[11]~FF  (.D(n2214), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[11]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[12]~FF  (.D(n2189), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[12]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[13]~FF  (.D(n2187), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[13]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[14]~FF  (.D(n2185), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[14]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[15]~FF  (.D(n2184), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[15]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[1]~FF  (.D(n946), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[2]~FF  (.D(n2179), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[3]~FF  (.D(n2177), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[4]~FF  (.D(n2175), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[5]~FF  (.D(n2173), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[6]~FF  (.D(n2171), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[7]~FF  (.D(n2169), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[8]~FF  (.D(n2167), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[9]~FF  (.D(n2165), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[10]~FF  (.D(n2163), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[11]~FF  (.D(n2161), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[12]~FF  (.D(n2159), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[13]~FF  (.D(n2157), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[14]~FF  (.D(n2155), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[15]~FF  (.D(n2154), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1162 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1161 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1160 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1159 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n885 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n884 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n883 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n882 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n881 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n880 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n879 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1179 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1178 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1177 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1176 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF  (.D(\u_scaler_gray/srcx_int[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF  (.D(\u_scaler_gray/srcx_int[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF  (.D(\u_scaler_gray/srcx_int[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF  (.D(\u_scaler_gray/srcx_int[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF  (.D(\u_scaler_gray/srcx_int[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF  (.D(\u_scaler_gray/srcx_int[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF  (.D(\u_scaler_gray/srcx_int[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1162 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1195 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1194 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1193 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1179 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1212 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1211 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1210 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/tvalid~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/tvalid )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/tvalid~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/tvalid~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/tvalid~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF  (.D(n910), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF  (.D(n2592), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF  (.D(n2590), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF  (.D(n2588), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF  (.D(n2586), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF  (.D(n2584), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF  (.D(n2582), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF  (.D(n2580), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF  (.D(n2578), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF  (.D(n2576), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF  (.D(n2574), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF  (.D(n2572), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF  (.D(n2570), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF  (.D(n2568), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF  (.D(n2555), 
           .CE(n197), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[1]~FF  (.D(\u_scaler_gray/n129 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[2]~FF  (.D(\u_scaler_gray/n128 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[3]~FF  (.D(\u_scaler_gray/n127 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[4]~FF  (.D(\u_scaler_gray/n126 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[5]~FF  (.D(\u_scaler_gray/n125 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[6]~FF  (.D(\u_scaler_gray/n124 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[7]~FF  (.D(\u_scaler_gray/n123 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[8]~FF  (.D(\u_scaler_gray/n122 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[9]~FF  (.D(\u_scaler_gray/n121 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[10]~FF  (.D(\u_scaler_gray/n120 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[11]~FF  (.D(\u_scaler_gray/n119 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[12]~FF  (.D(\u_scaler_gray/n118 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[12]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[13]~FF  (.D(\u_scaler_gray/n117 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[13]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[14]~FF  (.D(\u_scaler_gray/n116 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[14]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[15]~FF  (.D(\u_scaler_gray/n115 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[15]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n462 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ASIZE_0[2]~FF  (.D(1'b1), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(DdrCtrl_ALEN_0[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \DdrCtrl_ASIZE_0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ASIZE_0[2]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ASIZE_0[2]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ASIZE_0[2]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ASIZE_0[2]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_ASIZE_0[2]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ASIZE_0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF  (.D(n2152), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF  (.D(n2150), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF  (.D(n2148), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF  (.D(n2146), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF  (.D(n2142), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF  (.D(n2140), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF  (.D(n2138), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF  (.D(n2136), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF  (.D(n2134), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF  (.D(n2129), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF  (.D(n2125), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF  (.D(n2123), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF  (.D(n2119), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF  (.D(n2117), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF  (.D(n2115), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF  (.D(n2112), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF  (.D(n2110), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF  (.D(n1535), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF  (.D(n2107), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF  (.D(n2105), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF  (.D(n2102), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF  (.D(n2098), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF  (.D(n2096), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF  (.D(n2093), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF  (.D(n2091), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF  (.D(n2066), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF  (.D(n2064), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF  (.D(n2062), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF  (.D(n2060), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF  (.D(n2058), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF  (.D(n2056), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF  (.D(n2054), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF  (.D(n1783), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF  (.D(n1740), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF  (.D(n1706), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF  (.D(n1704), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF  (.D(n1702), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF  (.D(n1700), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF  (.D(n1698), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF  (.D(n1696), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF  (.D(n1694), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF  (.D(n1692), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF  (.D(n1690), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF  (.D(n1685), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__15140 (.I0(\u_axi4_ctrl/state[1] ), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(\u_axi4_ctrl/state[2] ), .O(DdrCtrl_AVALID_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__15140.LUTMASK = 16'h1414;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n335 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcx_fix[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n334 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcx_fix[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n333 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcx_fix[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n332 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n331 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n330 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n329 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n328 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n327 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n326 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n325 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[8]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n324 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n323 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n322 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n321 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[12]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n320 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[13]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n319 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[14]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n318 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[15]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n317 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n461 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n460 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n459 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n458 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n457 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n456 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n455 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n454 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n453 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n452 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n451 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n450 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n449 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n448 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n447 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n446 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n445 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n444 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n443 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[8]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n442 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n441 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n440 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n439 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[12]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n438 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[13]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n437 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[14]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n436 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[15]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n435 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF  (.D(\u_scaler_gray/destx[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF  (.D(\u_scaler_gray/destx[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF  (.D(n1537), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF  (.D(n1516), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF  (.D(n1514), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF  (.D(n1512), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF  (.D(n1510), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF  (.D(n1508), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF  (.D(n1506), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF  (.D(n1504), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF  (.D(n1502), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF  (.D(n1500), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF  (.D(n1498), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF  (.D(n1496), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF  (.D(n1494), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF  (.D(n1492), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF  (.D(n1490), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF  (.D(n1489), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(26)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcx_fix[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(26)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcx_fix[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(26)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcx_fix[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(26)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF  (.D(n1753), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF  (.D(n1918), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n344 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[0]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[0]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[0]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF  (.D(\u_scaler_gray/tvalid ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_GBUFCE CLKBUF__5 (.CE(1'b1), .I(jtag_inst1_TCK), .O(\jtag_inst1_TCK~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__5.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__4 (.CE(1'b1), .I(cmos_pclk), .O(\cmos_pclk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__4.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__3 (.CE(1'b1), .I(hdmi_clk2x_i), .O(\hdmi_clk2x_i~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__3.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__2 (.CE(1'b1), .I(hdmi_clk1x_i), .O(\hdmi_clk1x_i~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__2.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(tx_slowclk), .O(\tx_slowclk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF  (.D(n1115), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF  (.D(n1113), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF  (.D(n1109), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF  (.D(n1107), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF  (.D(n1105), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF  (.D(n1103), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF  (.D(n1101), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF  (.D(n1099), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF  (.D(n1097), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF  (.D(n1095), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF  (.D(n1093), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF  (.D(n1091), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF  (.D(n1089), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF  (.D(n1087), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF  (.D(n1085), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF  (.D(n1083), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF  (.D(n1081), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF  (.D(n1079), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF  (.D(n1077), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF  (.D(n1078), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF  (.D(n1075), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF  (.D(n1073), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF  (.D(n1071), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF  (.D(n1069), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF  (.D(n1067), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF  (.D(n1065), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF  (.D(n1063), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF  (.D(n1046), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF  (.D(n1044), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF  (.D(n1042), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF  (.D(n1040), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF  (.D(n1038), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF  (.D(n1036), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF  (.D(n1034), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF  (.D(n1032), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF  (.D(n1030), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF  (.D(n1028), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF  (.D(n1026), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF  (.D(n1024), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF  (.D(n1025), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF  (.D(n1012), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF  (.D(n1010), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF  (.D(n975), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF  (.D(n973), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF  (.D(n966), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF  (.D(n962), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF  (.D(n960), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF  (.D(n958), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF  (.D(n956), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF  (.D(n954), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF  (.D(n955), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n343 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n342 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n341 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n340 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n339 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n338 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n337 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n336 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n335 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[1]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[1]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[1]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[2]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[2]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[2]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[3]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[3]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[3]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[4]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[4]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[4]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[5]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[5]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[5]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[5]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[5]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[5]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[6]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[6]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[6]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[6]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[7]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[7]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[7]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[7]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tvalid_o~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(tvalid_o)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(70)
    defparam \tvalid_o~FF .CLK_POLARITY = 1'b1;
    defparam \tvalid_o~FF .CE_POLARITY = 1'b1;
    defparam \tvalid_o~FF .SR_POLARITY = 1'b1;
    defparam \tvalid_o~FF .D_POLARITY = 1'b1;
    defparam \tvalid_o~FF .SR_SYNC = 1'b1;
    defparam \tvalid_o~FF .SR_VALUE = 1'b0;
    defparam \tvalid_o~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(Axi_Clk), .O(\Axi_Clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_52/add_2/i2  (.I0(n3344), .I1(1'b1), 
            .CI(1'b0), .CO(n10608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(79)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_52/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_52/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_50/add_2/i2  (.I0(n3344), .I1(1'b1), 
            .CI(1'b0), .CO(n10607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_50/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_50/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__u_rgb2dvi/enc_2/sub_50/add_2/i1  (.I0(1'b0), .I1(1'b0), 
            .CI(n10606), .O(n3344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \AUX_ADD_CO__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_2/sub_50/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n10605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_79/add_2/i2  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n10604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(93)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_79/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_79/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n10603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n10602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n10601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n10599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n10598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n10597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n10596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20  (.I0(1'b0), 
            .I1(1'b0), .CI(n10595), .O(n1078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20  (.I0(1'b0), 
            .I1(1'b0), .CI(n10594), .O(n1025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21  (.I0(1'b0), 
            .I1(1'b0), .CI(n10593), .O(n955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n10592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \AUX_ADD_CI__u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n10591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[0]~FF  (.D(tvsync_o), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[0]~FF  (.D(lcd_vs), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_index[0]~FF  (.D(\u_axi4_ctrl/n317 ), .CE(\u_axi4_ctrl/equal_38/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(177)
    defparam \u_axi4_ctrl/wframe_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_index[0]~FF  (.D(\u_axi4_ctrl/n336 ), .CE(\u_axi4_ctrl/equal_47/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(197)
    defparam \u_axi4_ctrl/rframe_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/state[0]~FF  (.D(\u_axi4_ctrl/n389 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(268)
    defparam \u_axi4_ctrl/state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/state[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ATYPE_0~FF  (.D(1'b1), .CE(\u_axi4_ctrl/n405 ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/n1476 ), .Q(DdrCtrl_ATYPE_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(283)
    defparam \DdrCtrl_ATYPE_0~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ATYPE_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[0]~FF  (.D(\u_axi4_ctrl/wdata_cnt_dly[0] ), 
           .CE(\u_axi4_ctrl/n363 ), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), 
           .Q(\u_axi4_ctrl/wdata_cnt_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[1]~FF  (.D(\u_axi4_ctrl/n1544 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[0]~FF  (.D(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
           .CE(\u_axi4_ctrl/n379 ), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), 
           .Q(\u_axi4_ctrl/rdata_cnt_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wenb~FF  (.D(\u_axi4_ctrl/n379 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rfifo_wenb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(434)
    defparam \u_axi4_ctrl/rfifo_wenb~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[0]~FF  (.D(DdrCtrl_RDATA_0[0]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[1]~FF  (.D(\u_axi4_ctrl/wframe_vsync_dly[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[2]~FF  (.D(\u_axi4_ctrl/wframe_vsync_dly[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[3]~FF  (.D(\u_axi4_ctrl/wframe_vsync_dly[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[1]~FF  (.D(\u_axi4_ctrl/rframe_vsync_dly[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[2]~FF  (.D(\u_axi4_ctrl/rframe_vsync_dly[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[3]~FF  (.D(\u_axi4_ctrl/rframe_vsync_dly[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_index[1]~FF  (.D(\u_axi4_ctrl/n316 ), .CE(\u_axi4_ctrl/equal_38/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(177)
    defparam \u_axi4_ctrl/wframe_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF  (.D(n2340), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF  (.D(n2322), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wfifo_empty~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CE(ceg_net289), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/wfifo_empty )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1090)
    defparam \u_axi4_ctrl/wfifo_empty~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_empty~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_empty~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF  (.D(n755), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF  (.D(n753), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF  (.D(n751), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF  (.D(n749), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF  (.D(n747), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF  (.D(n726), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF  (.D(n722), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF  (.D(n717), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF  (.D(n696), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF  (.D(n693), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF  (.D(n2350), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF  (.D(n679), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF  (.D(n677), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF  (.D(n675), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF  (.D(n673), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF  (.D(n671), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF  (.D(n669), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF  (.D(n668), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_empty~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CE(ceg_net296), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/rfifo_empty )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1090)
    defparam \u_axi4_ctrl/rfifo_empty~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_empty~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_empty~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF  (.D(n2516), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF  (.D(n2519), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF  (.D(n564), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF  (.D(n562), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF  (.D(n560), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF  (.D(n558), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF  (.D(n556), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF  (.D(n555), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF  (.D(n2523), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF  (.D(n553), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF  (.D(n551), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF  (.D(n549), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF  (.D(n547), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF  (.D(n545), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF  (.D(n543), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF  (.D(n541), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF  (.D(n531), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF  (.D(n461), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF  (.D(n454), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF  (.D(n453), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32_q ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35  (.D(n10294), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_index[1]~FF  (.D(\u_axi4_ctrl/n335 ), .CE(\u_axi4_ctrl/equal_47/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(197)
    defparam \u_axi4_ctrl/rframe_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/state[1]~FF  (.D(\u_axi4_ctrl/n1612 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1619 ), .Q(\u_axi4_ctrl/state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(268)
    defparam \u_axi4_ctrl/state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/state[2]~FF  (.D(\u_axi4_ctrl/n387 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(268)
    defparam \u_axi4_ctrl/state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/state[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[10]~FF  (.D(\u_axi4_ctrl/awaddr[10] ), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[11]~FF  (.D(n1924), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[12]~FF  (.D(n928), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[13]~FF  (.D(n925), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[14]~FF  (.D(n921), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[15]~FF  (.D(n918), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[16]~FF  (.D(n914), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[17]~FF  (.D(n811), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[18]~FF  (.D(n809), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[19]~FF  (.D(n807), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[20]~FF  (.D(n805), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[21]~FF  (.D(n803), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[22]~FF  (.D(n801), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[23]~FF  (.D(n800), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[10]~FF  (.D(\u_axi4_ctrl/araddr[10] ), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[11]~FF  (.D(n2121), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[12]~FF  (.D(n798), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[13]~FF  (.D(n796), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[14]~FF  (.D(n794), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[15]~FF  (.D(n792), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[16]~FF  (.D(n790), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[17]~FF  (.D(n788), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[18]~FF  (.D(n786), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[19]~FF  (.D(n784), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[20]~FF  (.D(n782), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[21]~FF  (.D(n780), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[22]~FF  (.D(n778), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[23]~FF  (.D(n777), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[10]~FF  (.D(\u_axi4_ctrl/n697 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[10]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[10]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[10]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[11]~FF  (.D(\u_axi4_ctrl/n696 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[11]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[11]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[11]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[12]~FF  (.D(\u_axi4_ctrl/n695 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[12]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[12]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[12]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[13]~FF  (.D(\u_axi4_ctrl/n694 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[13]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[13]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[13]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[14]~FF  (.D(\u_axi4_ctrl/n693 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[14]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[14]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[14]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[15]~FF  (.D(\u_axi4_ctrl/n692 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[15]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[15]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[16]~FF  (.D(\u_axi4_ctrl/n691 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[16]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[16]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[16]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[17]~FF  (.D(\u_axi4_ctrl/n690 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[17]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[17]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[17]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[18]~FF  (.D(\u_axi4_ctrl/n689 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[18]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[18]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[18]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[19]~FF  (.D(\u_axi4_ctrl/n688 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[19]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[19]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[19]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[20]~FF  (.D(\u_axi4_ctrl/n687 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[20]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[20]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[20]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[21]~FF  (.D(\u_axi4_ctrl/n686 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[21]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[21]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[21]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[22]~FF  (.D(\u_axi4_ctrl/n685 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[22]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[22]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[22]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[23]~FF  (.D(\u_axi4_ctrl/n684 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[23]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[23]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[23]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[24]~FF  (.D(\u_axi4_ctrl/n683 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[24]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[24]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[24]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[25]~FF  (.D(\u_axi4_ctrl/n682 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[25]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[25]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[25]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[1]~FF  (.D(\u_axi4_ctrl/n1499 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[2]~FF  (.D(\u_axi4_ctrl/n1504 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[3]~FF  (.D(\u_axi4_ctrl/n1509 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[4]~FF  (.D(\u_axi4_ctrl/n1514 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[5]~FF  (.D(\u_axi4_ctrl/n1519 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[6]~FF  (.D(\u_axi4_ctrl/n1524 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[7]~FF  (.D(\u_axi4_ctrl/n1529 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[8]~FF  (.D(\u_axi4_ctrl/n1534 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[2]~FF  (.D(\u_axi4_ctrl/n1549 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[3]~FF  (.D(\u_axi4_ctrl/n1554 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[4]~FF  (.D(\u_axi4_ctrl/n1559 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[5]~FF  (.D(\u_axi4_ctrl/n1564 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[6]~FF  (.D(\u_axi4_ctrl/n1569 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[7]~FF  (.D(\u_axi4_ctrl/n1574 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[8]~FF  (.D(\u_axi4_ctrl/n1579 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[1]~FF  (.D(DdrCtrl_RDATA_0[1]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[2]~FF  (.D(DdrCtrl_RDATA_0[2]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[3]~FF  (.D(DdrCtrl_RDATA_0[3]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[4]~FF  (.D(DdrCtrl_RDATA_0[4]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[5]~FF  (.D(DdrCtrl_RDATA_0[5]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[6]~FF  (.D(DdrCtrl_RDATA_0[6]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[7]~FF  (.D(DdrCtrl_RDATA_0[7]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[8]~FF  (.D(DdrCtrl_RDATA_0[8]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[9]~FF  (.D(DdrCtrl_RDATA_0[9]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[10]~FF  (.D(DdrCtrl_RDATA_0[10]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[11]~FF  (.D(DdrCtrl_RDATA_0[11]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[12]~FF  (.D(DdrCtrl_RDATA_0[12]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[13]~FF  (.D(DdrCtrl_RDATA_0[13]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[14]~FF  (.D(DdrCtrl_RDATA_0[14]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[15]~FF  (.D(DdrCtrl_RDATA_0[15]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[16]~FF  (.D(DdrCtrl_RDATA_0[16]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[17]~FF  (.D(DdrCtrl_RDATA_0[17]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[18]~FF  (.D(DdrCtrl_RDATA_0[18]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[19]~FF  (.D(DdrCtrl_RDATA_0[19]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[20]~FF  (.D(DdrCtrl_RDATA_0[20]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[21]~FF  (.D(DdrCtrl_RDATA_0[21]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[22]~FF  (.D(DdrCtrl_RDATA_0[22]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[23]~FF  (.D(DdrCtrl_RDATA_0[23]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[24]~FF  (.D(DdrCtrl_RDATA_0[24]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[25]~FF  (.D(DdrCtrl_RDATA_0[25]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[26]~FF  (.D(DdrCtrl_RDATA_0[26]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[27]~FF  (.D(DdrCtrl_RDATA_0[27]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[28]~FF  (.D(DdrCtrl_RDATA_0[28]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[29]~FF  (.D(DdrCtrl_RDATA_0[29]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[30]~FF  (.D(DdrCtrl_RDATA_0[30]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[31]~FF  (.D(DdrCtrl_RDATA_0[31]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[32]~FF  (.D(DdrCtrl_RDATA_0[32]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[33]~FF  (.D(DdrCtrl_RDATA_0[33]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[34]~FF  (.D(DdrCtrl_RDATA_0[34]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[35]~FF  (.D(DdrCtrl_RDATA_0[35]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[36]~FF  (.D(DdrCtrl_RDATA_0[36]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[37]~FF  (.D(DdrCtrl_RDATA_0[37]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[38]~FF  (.D(DdrCtrl_RDATA_0[38]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[39]~FF  (.D(DdrCtrl_RDATA_0[39]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[40]~FF  (.D(DdrCtrl_RDATA_0[40]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[41]~FF  (.D(DdrCtrl_RDATA_0[41]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[42]~FF  (.D(DdrCtrl_RDATA_0[42]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[43]~FF  (.D(DdrCtrl_RDATA_0[43]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[44]~FF  (.D(DdrCtrl_RDATA_0[44]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[45]~FF  (.D(DdrCtrl_RDATA_0[45]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[46]~FF  (.D(DdrCtrl_RDATA_0[46]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[47]~FF  (.D(DdrCtrl_RDATA_0[47]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[48]~FF  (.D(DdrCtrl_RDATA_0[48]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[49]~FF  (.D(DdrCtrl_RDATA_0[49]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[50]~FF  (.D(DdrCtrl_RDATA_0[50]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[51]~FF  (.D(DdrCtrl_RDATA_0[51]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[52]~FF  (.D(DdrCtrl_RDATA_0[52]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[53]~FF  (.D(DdrCtrl_RDATA_0[53]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[54]~FF  (.D(DdrCtrl_RDATA_0[54]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[55]~FF  (.D(DdrCtrl_RDATA_0[55]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[56]~FF  (.D(DdrCtrl_RDATA_0[56]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[57]~FF  (.D(DdrCtrl_RDATA_0[57]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[58]~FF  (.D(DdrCtrl_RDATA_0[58]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[59]~FF  (.D(DdrCtrl_RDATA_0[59]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[60]~FF  (.D(DdrCtrl_RDATA_0[60]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[61]~FF  (.D(DdrCtrl_RDATA_0[61]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[62]~FF  (.D(DdrCtrl_RDATA_0[62]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[63]~FF  (.D(DdrCtrl_RDATA_0[63]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[64]~FF  (.D(DdrCtrl_RDATA_0[64]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[65]~FF  (.D(DdrCtrl_RDATA_0[65]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[66]~FF  (.D(DdrCtrl_RDATA_0[66]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[67]~FF  (.D(DdrCtrl_RDATA_0[67]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[68]~FF  (.D(DdrCtrl_RDATA_0[68]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[69]~FF  (.D(DdrCtrl_RDATA_0[69]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[70]~FF  (.D(DdrCtrl_RDATA_0[70]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[71]~FF  (.D(DdrCtrl_RDATA_0[71]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[72]~FF  (.D(DdrCtrl_RDATA_0[72]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[73]~FF  (.D(DdrCtrl_RDATA_0[73]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[74]~FF  (.D(DdrCtrl_RDATA_0[74]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[75]~FF  (.D(DdrCtrl_RDATA_0[75]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[76]~FF  (.D(DdrCtrl_RDATA_0[76]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[77]~FF  (.D(DdrCtrl_RDATA_0[77]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[78]~FF  (.D(DdrCtrl_RDATA_0[78]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[79]~FF  (.D(DdrCtrl_RDATA_0[79]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[80]~FF  (.D(DdrCtrl_RDATA_0[80]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[81]~FF  (.D(DdrCtrl_RDATA_0[81]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[82]~FF  (.D(DdrCtrl_RDATA_0[82]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[83]~FF  (.D(DdrCtrl_RDATA_0[83]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[84]~FF  (.D(DdrCtrl_RDATA_0[84]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[85]~FF  (.D(DdrCtrl_RDATA_0[85]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[86]~FF  (.D(DdrCtrl_RDATA_0[86]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[87]~FF  (.D(DdrCtrl_RDATA_0[87]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[88]~FF  (.D(DdrCtrl_RDATA_0[88]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[89]~FF  (.D(DdrCtrl_RDATA_0[89]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[90]~FF  (.D(DdrCtrl_RDATA_0[90]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[91]~FF  (.D(DdrCtrl_RDATA_0[91]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[92]~FF  (.D(DdrCtrl_RDATA_0[92]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[93]~FF  (.D(DdrCtrl_RDATA_0[93]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[94]~FF  (.D(DdrCtrl_RDATA_0[94]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[95]~FF  (.D(DdrCtrl_RDATA_0[95]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[96]~FF  (.D(DdrCtrl_RDATA_0[96]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[97]~FF  (.D(DdrCtrl_RDATA_0[97]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[98]~FF  (.D(DdrCtrl_RDATA_0[98]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[99]~FF  (.D(DdrCtrl_RDATA_0[99]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[100]~FF  (.D(DdrCtrl_RDATA_0[100]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[101]~FF  (.D(DdrCtrl_RDATA_0[101]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[102]~FF  (.D(DdrCtrl_RDATA_0[102]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[103]~FF  (.D(DdrCtrl_RDATA_0[103]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[104]~FF  (.D(DdrCtrl_RDATA_0[104]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[105]~FF  (.D(DdrCtrl_RDATA_0[105]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[106]~FF  (.D(DdrCtrl_RDATA_0[106]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[107]~FF  (.D(DdrCtrl_RDATA_0[107]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[108]~FF  (.D(DdrCtrl_RDATA_0[108]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[109]~FF  (.D(DdrCtrl_RDATA_0[109]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[110]~FF  (.D(DdrCtrl_RDATA_0[110]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[111]~FF  (.D(DdrCtrl_RDATA_0[111]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[112]~FF  (.D(DdrCtrl_RDATA_0[112]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[113]~FF  (.D(DdrCtrl_RDATA_0[113]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[114]~FF  (.D(DdrCtrl_RDATA_0[114]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[115]~FF  (.D(DdrCtrl_RDATA_0[115]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[116]~FF  (.D(DdrCtrl_RDATA_0[116]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[117]~FF  (.D(DdrCtrl_RDATA_0[117]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[118]~FF  (.D(DdrCtrl_RDATA_0[118]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[119]~FF  (.D(DdrCtrl_RDATA_0[119]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[120]~FF  (.D(DdrCtrl_RDATA_0[120]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[121]~FF  (.D(DdrCtrl_RDATA_0[121]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[122]~FF  (.D(DdrCtrl_RDATA_0[122]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[123]~FF  (.D(DdrCtrl_RDATA_0[123]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[124]~FF  (.D(DdrCtrl_RDATA_0[124]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[125]~FF  (.D(DdrCtrl_RDATA_0[125]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[126]~FF  (.D(DdrCtrl_RDATA_0[126]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[127]~FF  (.D(DdrCtrl_RDATA_0[127]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[0]~FF  (.D(\u_lcd_driver/n83 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_hs~FF  (.D(\u_lcd_driver/n35 ), .CE(r_hdmi_rst_n), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(lcd_hs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \lcd_hs~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_hs~FF .CE_POLARITY = 1'b1;
    defparam \lcd_hs~FF .SR_POLARITY = 1'b1;
    defparam \lcd_hs~FF .D_POLARITY = 1'b0;
    defparam \lcd_hs~FF .SR_SYNC = 1'b1;
    defparam \lcd_hs~FF .SR_VALUE = 1'b0;
    defparam \lcd_hs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_vs~FF  (.D(\u_lcd_driver/n97 ), .CE(r_hdmi_rst_n), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(lcd_vs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \lcd_vs~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_vs~FF .CE_POLARITY = 1'b1;
    defparam \lcd_vs~FF .SR_POLARITY = 1'b1;
    defparam \lcd_vs~FF .D_POLARITY = 1'b0;
    defparam \lcd_vs~FF .SR_SYNC = 1'b1;
    defparam \lcd_vs~FF .SR_VALUE = 1'b0;
    defparam \lcd_vs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_de~FF  (.D(\u_lcd_driver/n125 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(lcd_de)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \lcd_de~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_de~FF .CE_POLARITY = 1'b1;
    defparam \lcd_de~FF .SR_POLARITY = 1'b1;
    defparam \lcd_de~FF .D_POLARITY = 1'b1;
    defparam \lcd_de~FF .SR_SYNC = 1'b1;
    defparam \lcd_de~FF .SR_VALUE = 1'b0;
    defparam \lcd_de~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_dv~FF  (.D(\u_lcd_driver/n133 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_dv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_dv~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[0]~FF  (.D(\u_lcd_driver/n34 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[1]~FF  (.D(\u_lcd_driver/n82 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[2]~FF  (.D(\u_lcd_driver/n81 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[3]~FF  (.D(\u_lcd_driver/n80 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[4]~FF  (.D(\u_lcd_driver/n79 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[5]~FF  (.D(\u_lcd_driver/n78 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[6]~FF  (.D(\u_lcd_driver/n77 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[7]~FF  (.D(\u_lcd_driver/n76 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[8]~FF  (.D(\u_lcd_driver/n75 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[9]~FF  (.D(\u_lcd_driver/n74 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[10]~FF  (.D(\u_lcd_driver/n73 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[11]~FF  (.D(\u_lcd_driver/n72 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__15141 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/wdata_cnt_dly[3] ), 
            .O(n10069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15141.LUTMASK = 16'h8000;
    EFX_FF \u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36  (.D(n10292), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true", INIT_VALUE=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32 .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32 .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32 .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32 .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32 .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32 .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37  (.D(n10290), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37 .D_POLARITY = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[1]~FF  (.D(\u_lcd_driver/n33 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[2]~FF  (.D(\u_lcd_driver/n32 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[3]~FF  (.D(\u_lcd_driver/n31 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[4]~FF  (.D(\u_lcd_driver/n30 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[5]~FF  (.D(\u_lcd_driver/n29 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[6]~FF  (.D(\u_lcd_driver/n28 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[7]~FF  (.D(\u_lcd_driver/n27 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[8]~FF  (.D(\u_lcd_driver/n26 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[9]~FF  (.D(\u_lcd_driver/n25 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[10]~FF  (.D(\u_lcd_driver/n24 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[11]~FF  (.D(\u_lcd_driver/n23 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[0]~FF  (.D(\u_rgb2dvi/enc_0/n866 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[0]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[0]~FF  (.D(n3203), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_0/acc[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[1]~FF  (.D(\u_rgb2dvi/enc_0/n768 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[1]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[1]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[1]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[1]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[1]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[1]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[2]~FF  (.D(\u_rgb2dvi/enc_0/n774 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[2]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[2]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[2]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[2]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[2]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[3]~FF  (.D(\u_rgb2dvi/enc_0/n780 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[3]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[3]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[3]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[3]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[3]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[3]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[4]~FF  (.D(\u_rgb2dvi/enc_0/n786 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[4]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[4]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[5]~FF  (.D(\u_rgb2dvi/enc_0/n792 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[5]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[5]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[5]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[5]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[5]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[5]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[6]~FF  (.D(\u_rgb2dvi/enc_0/n798 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[6]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[6]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[6]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[6]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[6]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[6]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[7]~FF  (.D(\u_rgb2dvi/enc_0/n804 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[7]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[7]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[7]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[7]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[7]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[7]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[8]~FF  (.D(\u_rgb2dvi/enc_0/n810 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[8]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[8]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[9]~FF  (.D(\u_rgb2dvi/enc_0/n816 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[9]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[9]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[1]~FF  (.D(n385), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_0/acc[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[2]~FF  (.D(n383), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_0/acc[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[3]~FF  (.D(n381), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_0/acc[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[4]~FF  (.D(n380), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_0/acc[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[0]~FF  (.D(\u_rgb2dvi/enc_1/q_out[0] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[0]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[0]~FF  (.D(n3282), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_1/acc[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[1]~FF  (.D(\u_rgb2dvi/enc_1/q_out[1] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[1]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[1]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[1]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[1]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[1]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[2]~FF  (.D(\u_rgb2dvi/enc_1/q_out[2] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[2]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[2]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[2]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[2]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[2]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[3]~FF  (.D(\u_rgb2dvi/enc_1/q_out[3] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[3]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[3]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[3]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[3]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[3]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[4]~FF  (.D(\u_rgb2dvi/enc_1/q_out[4] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[4]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[4]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[4]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[4]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[4]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[5]~FF  (.D(\u_rgb2dvi/enc_1/q_out[5] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[5]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[5]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[5]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[5]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[5]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[6]~FF  (.D(\u_rgb2dvi/enc_1/q_out[6] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[6]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[6]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[6]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[6]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[6]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[7]~FF  (.D(\u_rgb2dvi/enc_1/q_out[7] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[7]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[7]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[7]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[7]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[7]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[8]~FF  (.D(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q_pinv ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[8]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[9]~FF  (.D(\u_rgb2dvi/enc_1/q_out[9] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[9]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[9]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[9]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[9]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[9]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[1]~FF  (.D(n359), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_1/acc[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[2]~FF  (.D(n357), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_1/acc[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[3]~FF  (.D(n355), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_1/acc[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[4]~FF  (.D(n354), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_1/acc[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[0]~FF  (.D(\u_rgb2dvi/enc_2/q_out[0] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[0]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[0]~FF  (.D(n3339), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_2/acc[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[1]~FF  (.D(\u_rgb2dvi/enc_2/q_out[1] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[1]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[1]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[1]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[1]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[1]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[2]~FF  (.D(\u_rgb2dvi/enc_2/q_out[2] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[2]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[2]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[2]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[2]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[2]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[3]~FF  (.D(\u_rgb2dvi/enc_2/q_out[3] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[3]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[3]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[3]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[3]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[3]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[4]~FF  (.D(\u_rgb2dvi/enc_2/q_out[4] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[4]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[4]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[4]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[4]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[4]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[5]~FF  (.D(\u_rgb2dvi/enc_2/q_out[5] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[5]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[5]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[5]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[5]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[5]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[6]~FF  (.D(\u_rgb2dvi/enc_2/q_out[6] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[6]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[6]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[6]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[6]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[6]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[7]~FF  (.D(\u_rgb2dvi/enc_2/q_out[7] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[7]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[7]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[7]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[7]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[7]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[9]~FF  (.D(\u_rgb2dvi/enc_2/q_out[9] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[9]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[9]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[9]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[9]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[9]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[1]~FF  (.D(n350), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_2/acc[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[2]~FF  (.D(n348), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_2/acc[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[3]~FF  (.D(n346), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_2/acc[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[4]~FF  (.D(n345), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_2/acc[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_txc_o[1]~FF  (.D(\r_hdmi_txc_o[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(hdmi_txc_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_txc_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_txc_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_txc_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_txc_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_txc_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_txc_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_txc_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_txc_o[9]~FF  (.D(rc_hdmi_tx), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(\r_hdmi_txc_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_txc_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .SR_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_txc_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[1]~FF  (.D(n591), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx0_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[2]~FF  (.D(n590), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx0_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[3]~FF  (.D(n589), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx0_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[4]~FF  (.D(n588), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx0_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[5]~FF  (.D(\w_hdmi_txd0[5] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx0_o[5]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[5]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[5]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[5]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[5]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[5]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[6]~FF  (.D(\w_hdmi_txd0[6] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx0_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[6]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[6]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[6]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[7]~FF  (.D(\w_hdmi_txd0[7] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx0_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[7]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[8]~FF  (.D(\w_hdmi_txd0[8] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx0_o[8]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[8]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[8]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[8]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[8]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[8]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[9]~FF  (.D(\w_hdmi_txd0[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx0_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[9]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[1]~FF  (.D(n602_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx1_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[2]~FF  (.D(n601_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx1_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[3]~FF  (.D(n600_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx1_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[4]~FF  (.D(n599_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx1_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[5]~FF  (.D(\w_hdmi_txd1[5] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx1_o[5]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[5]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[5]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[5]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[5]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[5]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[6]~FF  (.D(\w_hdmi_txd1[6] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx1_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[6]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[6]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[6]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[7]~FF  (.D(\w_hdmi_txd1[7] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx1_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[7]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[8]~FF  (.D(\w_hdmi_txd1[8] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx1_o[8]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[8]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[8]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[8]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[8]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[8]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[9]~FF  (.D(\w_hdmi_txd1[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx1_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[9]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[1]~FF  (.D(n613), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx2_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[2]~FF  (.D(n612), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx2_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[3]~FF  (.D(n611), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx2_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[4]~FF  (.D(n610), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx2_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[5]~FF  (.D(\w_hdmi_txd2[5] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx2_o[5]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[5]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[5]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[5]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[5]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[5]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[6]~FF  (.D(\w_hdmi_txd2[6] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx2_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[6]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[6]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[6]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[7]~FF  (.D(\w_hdmi_txd2[7] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx2_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[7]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[9]~FF  (.D(\w_hdmi_txd2[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx2_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[9]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[1]~FF  (.D(n4988), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[2]~FF  (.D(n4986), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[3]~FF  (.D(n4984), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[4]~FF  (.D(n3441), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[5]~FF  (.D(n3439), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[6]~FF  (.D(n3437), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[7]~FF  (.D(n3436), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig~FF  (.D(\edb_top_inst/la0/n1317 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_run_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig_imdt~FF  (.D(\edb_top_inst/la0/n1318 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig_imdt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_stop_trig~FF  (.D(\edb_top_inst/la0/n1319 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_stop_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_stop_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[0]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[0]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_soft_reset_in~FF  (.D(\edb_top_inst/la0/n1942 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_soft_reset_in )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3643)
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[0]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[0] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3672)
    defparam \edb_top_inst/la0/opcode[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[0]~FF  (.D(\edb_top_inst/la0/n2166 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[0]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[0] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[0]~FF  (.D(\edb_top_inst/la0/n2443 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[0]~FF  (.D(\edb_top_inst/la0/module_next_state[0] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3754)
    defparam \edb_top_inst/la0/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn_p1~FF  (.D(1'b1), .CE(1'b1), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/n2730 ), .Q(\edb_top_inst/la0/la_resetn_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4064)
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n2743 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4183)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n2743 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4183)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn~FF  (.D(\edb_top_inst/la0/la_resetn_p1 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/n2730 ), 
           .Q(\edb_top_inst/la0/la_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4064)
    defparam \edb_top_inst/la0/la_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF  (.D(lcd_vs), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4091)
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n2743 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4183)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF  (.D(lcd_de), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4091)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3576 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4183)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3576 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4183)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF  (.D(\lcd_data[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4091)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4465 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4183)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4480 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4678 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4400)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[0]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[0]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[32]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[33]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[34]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[35]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[36]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[37]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[38]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[39]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[40]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[41]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[42]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[43]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[44]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[45]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[46]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[47]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[48]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[49]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[50]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[51]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[52]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[53]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[54]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[55]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[56]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[57]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[58]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[59]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[60]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[61]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[62]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[63]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1373 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3616)
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[1]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[2]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[3]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[4]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[5]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[6]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[7]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[8]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[9]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[10]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[11]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[12]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[13]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[14]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[15]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[16]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[1]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[2]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[3]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[4]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1890 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3628)
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[1]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[1] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[2]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[2] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[3]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[3] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[4]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[4] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[5]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[5] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[6]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[6] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[7]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[7] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[8]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[8] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[9]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[9] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[10]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[10] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[11]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[11] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[12]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[12] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[13]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[13] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[14]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[14] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[15]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[15] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[16]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[16] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[17]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[17] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[18]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[18] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[19]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[19] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[20]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[20] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[21]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[21] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[22]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[22] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[23]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[23] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[24]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[24] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[25]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[25] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[26]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[26] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/address_counter[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3672)
    defparam \edb_top_inst/la0/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3672)
    defparam \edb_top_inst/la0/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3672)
    defparam \edb_top_inst/la0/opcode[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[1]~FF  (.D(\edb_top_inst/la0/n2165 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[2]~FF  (.D(\edb_top_inst/la0/n2164 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[3]~FF  (.D(\edb_top_inst/la0/n2163 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[4]~FF  (.D(\edb_top_inst/la0/n2162 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[5]~FF  (.D(\edb_top_inst/la0/n2161 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[1]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[1] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[2]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[2] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[3]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[3] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[4]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[4] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[5]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[5] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[6]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[6] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[7]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[7] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[8]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[8] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[9]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[9] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[10]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[10] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[11]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[11] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[12]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[12] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[13]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[13] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[14]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[14] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[15]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[15] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3699)
    defparam \edb_top_inst/la0/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[1]~FF  (.D(\edb_top_inst/la0/n2442 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[2]~FF  (.D(\edb_top_inst/la0/n2441 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[3]~FF  (.D(\edb_top_inst/la0/n2440 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[4]~FF  (.D(\edb_top_inst/la0/n2439 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[5]~FF  (.D(\edb_top_inst/la0/n2438 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[6]~FF  (.D(\edb_top_inst/la0/n2437 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[7]~FF  (.D(\edb_top_inst/la0/n2436 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[8]~FF  (.D(\edb_top_inst/la0/n2435 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[9]~FF  (.D(\edb_top_inst/la0/n2434 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[10]~FF  (.D(\edb_top_inst/la0/n2433 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[11]~FF  (.D(\edb_top_inst/la0/n2432 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[12]~FF  (.D(\edb_top_inst/la0/n2431 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[13]~FF  (.D(\edb_top_inst/la0/n2430 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[14]~FF  (.D(\edb_top_inst/la0/n2429 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[15]~FF  (.D(\edb_top_inst/la0/n2428 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[16]~FF  (.D(\edb_top_inst/la0/n2427 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[17]~FF  (.D(\edb_top_inst/la0/n2426 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[18]~FF  (.D(\edb_top_inst/la0/n2425 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[19]~FF  (.D(\edb_top_inst/la0/n2424 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[20]~FF  (.D(\edb_top_inst/la0/n2423 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[21]~FF  (.D(\edb_top_inst/la0/n2422 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[22]~FF  (.D(\edb_top_inst/la0/n2421 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[23]~FF  (.D(\edb_top_inst/la0/n2420 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[24]~FF  (.D(\edb_top_inst/la0/n2419 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[25]~FF  (.D(\edb_top_inst/la0/n2418 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[26]~FF  (.D(\edb_top_inst/la0/n2417 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[27]~FF  (.D(\edb_top_inst/la0/n2416 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[28]~FF  (.D(\edb_top_inst/la0/n2415 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[29]~FF  (.D(\edb_top_inst/la0/n2414 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[30]~FF  (.D(\edb_top_inst/la0/n2413 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[31]~FF  (.D(\edb_top_inst/la0/n2412 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[32]~FF  (.D(\edb_top_inst/la0/n2411 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[33]~FF  (.D(\edb_top_inst/la0/n2410 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[34]~FF  (.D(\edb_top_inst/la0/n2409 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[35]~FF  (.D(\edb_top_inst/la0/n2408 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[36]~FF  (.D(\edb_top_inst/la0/n2407 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[37]~FF  (.D(\edb_top_inst/la0/n2406 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[38]~FF  (.D(\edb_top_inst/la0/n2405 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[39]~FF  (.D(\edb_top_inst/la0/n2404 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[40]~FF  (.D(\edb_top_inst/la0/n2403 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[41]~FF  (.D(\edb_top_inst/la0/n2402 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[42]~FF  (.D(\edb_top_inst/la0/n2401 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[43]~FF  (.D(\edb_top_inst/la0/n2400 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[44]~FF  (.D(\edb_top_inst/la0/n2399 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[45]~FF  (.D(\edb_top_inst/la0/n2398 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[46]~FF  (.D(\edb_top_inst/la0/n2397 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[47]~FF  (.D(\edb_top_inst/la0/n2396 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[48]~FF  (.D(\edb_top_inst/la0/n2395 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[49]~FF  (.D(\edb_top_inst/la0/n2394 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[50]~FF  (.D(\edb_top_inst/la0/n2393 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[51]~FF  (.D(\edb_top_inst/la0/n2392 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[52]~FF  (.D(\edb_top_inst/la0/n2391 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[53]~FF  (.D(\edb_top_inst/la0/n2390 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[54]~FF  (.D(\edb_top_inst/la0/n2389 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[55]~FF  (.D(\edb_top_inst/la0/n2388 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[56]~FF  (.D(\edb_top_inst/la0/n2387 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[57]~FF  (.D(\edb_top_inst/la0/n2386 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[58]~FF  (.D(\edb_top_inst/la0/n2385 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[59]~FF  (.D(\edb_top_inst/la0/n2384 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[60]~FF  (.D(\edb_top_inst/la0/n2383 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[61]~FF  (.D(\edb_top_inst/la0/n2382 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[62]~FF  (.D(\edb_top_inst/la0/n2381 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[63]~FF  (.D(\edb_top_inst/la0/n2380 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3712)
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[1]~FF  (.D(\edb_top_inst/la0/module_next_state[1] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3754)
    defparam \edb_top_inst/la0/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[2]~FF  (.D(\edb_top_inst/la0/module_next_state[2] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3754)
    defparam \edb_top_inst/la0/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[3]~FF  (.D(\edb_top_inst/la0/module_next_state[3] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3754)
    defparam \edb_top_inst/la0/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[0]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n150 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[1]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n149 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[2]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n148 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[3]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n147 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[4]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n146 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[5]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n145 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[6]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n144 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[7]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n143 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[8]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n142 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[9]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n141 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[10]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n140 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[11]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n139 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[12]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n138 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[13]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n137 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[14]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n136 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[15]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n135 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[16]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n134 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[17]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n133 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[18]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n132 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[19]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n131 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[20]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n130 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[21]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n129 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[22]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n128 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[23]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n127 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[24]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n126 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[25]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n125 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[26]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n124 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[27]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n123 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[28]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n122 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[29]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n121 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[30]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n120 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[31]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n119 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(244)
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n19 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5482)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n3576 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4183)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF  (.D(\lcd_data[1] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4091)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF  (.D(\lcd_data[2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4091)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF  (.D(\lcd_data[3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4091)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF  (.D(\lcd_data[4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4091)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF  (.D(\lcd_data[5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4091)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF  (.D(\lcd_data[6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4091)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF  (.D(\lcd_data[7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4091)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5482)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n19 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5543)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5482)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4465 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4183)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4465 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4183)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4480 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4480 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n4480 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n4480 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n4480 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n4480 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n4480 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4199)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4678 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4678 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n4678 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n4678 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n4678 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n4678 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n4678 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4215)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n21 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n20 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n19 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5594)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/tu_trigger~FF  (.D(\edb_top_inst/la0/trigger_tu/n35 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/tu_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5724)
    defparam \edb_top_inst/la0/tu_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[2]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[3]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[4]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[5]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[6]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[7]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[8]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[9]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4388)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[1] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4400)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4400)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[3]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4400)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[4]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4400)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4400)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4400)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[7]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4400)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[8]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[8] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4400)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[9]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[9] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4400)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5210)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5010)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF  (.D(\edb_top_inst/la0/la_run_trig_imdt ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5010)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5010)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/str_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5231)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5246)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5246)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5246)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5256)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5269)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5269)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5269)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[0] ), 
           .CE(\edb_top_inst/ceg_net351 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5393)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1236 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/n7224 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5210)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5210)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[1] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5210)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF  (.D(\edb_top_inst/la0/la_run_trig ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5010)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/biu_ready~FF  (.D(\edb_top_inst/la0/la_biu_inst/n350 ), 
           .CE(\edb_top_inst/ceg_net348 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/biu_ready )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5281)
    defparam \edb_top_inst/la0/biu_ready~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF  (.D(\edb_top_inst/la0/address_counter[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF  (.D(\edb_top_inst/la0/address_counter[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF  (.D(\edb_top_inst/la0/address_counter[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF  (.D(\edb_top_inst/la0/address_counter[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF  (.D(\edb_top_inst/la0/address_counter[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF  (.D(\edb_top_inst/la0/address_counter[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF  (.D(\edb_top_inst/la0/address_counter[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF  (.D(\edb_top_inst/la0/address_counter[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF  (.D(\edb_top_inst/la0/address_counter[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF  (.D(\edb_top_inst/la0/address_counter[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF  (.D(\edb_top_inst/la0/address_counter[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF  (.D(\edb_top_inst/la0/address_counter[26] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n350 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5291)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[1] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[2] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[3] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[4] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[5] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[6] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[7] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[8] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[9] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[10] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1251 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_resetn ), .Q(\edb_top_inst/la0/data_from_biu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5300)
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] ), 
           .CE(\edb_top_inst/ceg_net351 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(5393)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[0]~FF  (.D(\edb_top_inst/la0/la_sample_cnt[0] ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_push ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/n1993 ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF  (.D(\edb_top_inst/n297 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF  (.D(\edb_top_inst/n765 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF  (.D(\edb_top_inst/n763 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF  (.D(\edb_top_inst/n761 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF  (.D(\edb_top_inst/n759 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF  (.D(\edb_top_inst/n757 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF  (.D(\edb_top_inst/n755 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF  (.D(\edb_top_inst/n753 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF  (.D(\edb_top_inst/n751 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF  (.D(\edb_top_inst/n749 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF  (.D(\edb_top_inst/n748 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF  (.D(\edb_top_inst/n426 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF  (.D(\edb_top_inst/n746 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF  (.D(\edb_top_inst/n744 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF  (.D(\edb_top_inst/n742 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF  (.D(\edb_top_inst/n740 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF  (.D(\edb_top_inst/n738 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF  (.D(\edb_top_inst/n736 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF  (.D(\edb_top_inst/n734 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF  (.D(\edb_top_inst/n732 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF  (.D(\edb_top_inst/n730 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF  (.D(\edb_top_inst/n727 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1993 ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF  (.D(\edb_top_inst/n428 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF  (.D(\edb_top_inst/n695 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF  (.D(\edb_top_inst/n693 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF  (.D(\edb_top_inst/n691 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF  (.D(\edb_top_inst/n689 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF  (.D(\edb_top_inst/n687 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF  (.D(\edb_top_inst/n685 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF  (.D(\edb_top_inst/n683 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF  (.D(\edb_top_inst/n681 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF  (.D(\edb_top_inst/n679 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF  (.D(\edb_top_inst/n677 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\tx_slowclk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[1]~FF  (.D(\edb_top_inst/n434 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[2]~FF  (.D(\edb_top_inst/n630 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[3]~FF  (.D(\edb_top_inst/n628 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[4]~FF  (.D(\edb_top_inst/n626 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[5]~FF  (.D(\edb_top_inst/n624 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[6]~FF  (.D(\edb_top_inst/n622 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[7]~FF  (.D(\edb_top_inst/n620 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[8]~FF  (.D(\edb_top_inst/n618 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[9]~FF  (.D(\edb_top_inst/n616 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[10]~FF  (.D(\edb_top_inst/n614 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[11]~FF  (.D(\edb_top_inst/n612 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[12]~FF  (.D(\edb_top_inst/n590 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4640)
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[1] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[8] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[9] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4709)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4531)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF  (.D(\edb_top_inst/n432 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF  (.D(\edb_top_inst/n651 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF  (.D(\edb_top_inst/n649 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF  (.D(\edb_top_inst/n647 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF  (.D(\edb_top_inst/n645 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF  (.D(\edb_top_inst/n643 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF  (.D(\edb_top_inst/n641 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF  (.D(\edb_top_inst/n639 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF  (.D(\edb_top_inst/n637 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF  (.D(\edb_top_inst/n635 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF  (.D(\edb_top_inst/n633 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF  (.D(\edb_top_inst/n632 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\tx_slowclk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4626)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[1]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[2]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[3]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[4]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[5]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[6]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[7]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[8]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[9]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[10]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[11]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[12]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3557)
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[1]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[2]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[3]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[4]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[5]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[6]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[7]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[8]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[9]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[10]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[11]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[12]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[13]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[14]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[15]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[16]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n6737 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3606)
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(315)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[0]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(315)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(315)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(315)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[1]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[2]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[3]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[4]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[5]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[6]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[7]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[8]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[9]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[10]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[11]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[12]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[13]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[14]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[15]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[16]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[17]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[18]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[19]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[20]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[21]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[22]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[23]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[24]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[25]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[26]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[27]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[28]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[29]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[30]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[31]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[32]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[33]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[34]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[35]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[36]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[37]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[38]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[39]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[40]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[41]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[42]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[43]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[44]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[45]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[46]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[47]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[48]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[49]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[50]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[51]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[52]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[53]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[54]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[55]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[56]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[57]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[58]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[59]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[60]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[61]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[62]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[63]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[64]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[65]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[66]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[67]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[68]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[69]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[70]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[71]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[72]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[73]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[74]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[75]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[76]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[77]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[78]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[79]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[80]~FF  (.D(\edb_top_inst/edb_user_dr[81] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[81]~FF  (.D(jtag_inst1_TDI), .CE(\edb_top_inst/debug_hub_inst/n95 ), 
           .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(308)
    defparam \edb_top_inst/edb_user_dr[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] ), 
            .I1(1'b0), .CI(n10591), .O(n186), .CO(n187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i2  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0] ), .CI(1'b0), 
            .O(n205), .CO(n206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i2 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i2  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] ), .CI(1'b0), 
            .O(n228), .CO(n229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i2 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i2  (.I0(\i2c_config_index[1] ), 
            .I1(\i2c_config_index[0] ), .CI(1'b0), .O(n231), .CO(n232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i2 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i5  (.I0(\u_rgb2dvi/enc_2/acc[4] ), .I1(n5371), 
            .CI(n347), .O(n345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i4  (.I0(\u_rgb2dvi/enc_2/acc[3] ), .I1(n5374), 
            .CI(n349), .O(n346), .CO(n347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i3  (.I0(\u_rgb2dvi/enc_2/acc[2] ), .I1(n5377), 
            .CI(n351), .O(n348), .CO(n349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i2  (.I0(\u_rgb2dvi/enc_2/acc[1] ), .I1(n5380), 
            .CI(n3340), .O(n350), .CO(n351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_75/i4  (.I0(n367), .I1(1'b0), .CI(n389), 
            .O(n352), .CO(n353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_2/add_75/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_75/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i5  (.I0(\u_rgb2dvi/enc_1/acc[4] ), .I1(n5385), 
            .CI(n356), .O(n354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i4  (.I0(\u_rgb2dvi/enc_1/acc[3] ), .I1(n5388), 
            .CI(n358), .O(n355), .CO(n356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i3  (.I0(\u_rgb2dvi/enc_1/acc[2] ), .I1(n5391), 
            .CI(n360), .O(n357), .CO(n358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i2  (.I0(\u_rgb2dvi/enc_1/acc[1] ), .I1(n5394), 
            .CI(n3283), .O(n359), .CO(n360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i5  (.I0(n373), .I1(1'b1), .CI(n363), 
            .O(n361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i4  (.I0(n374), .I1(1'b1), .CI(n365), 
            .O(n362), .CO(n363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i3  (.I0(n376), .I1(1'b1), .CI(n3218), 
            .O(n364), .CO(n365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i5  (.I0(1'b0), .I1(1'b1), .CI(n368), 
            .O(n366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i4  (.I0(n5403), .I1(n5413), .CI(n370), 
            .O(n367), .CO(n368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i3  (.I0(n5417), .I1(n5416), .CI(n372), 
            .O(n369), .CO(n370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i3 .I0_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i2  (.I0(n5420), .I1(n5410), .CI(n10608), 
            .O(n371), .CO(n372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i2 .I0_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i5  (.I0(1'b0), .I1(1'b1), .CI(n375), 
            .O(n373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i4  (.I0(n5413), .I1(n5403), .CI(n377), 
            .O(n374), .CO(n375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i3  (.I0(n5416), .I1(n5417), .CI(n379), 
            .O(n376), .CO(n377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i2  (.I0(n5410), .I1(n5420), .CI(n10607), 
            .O(n378), .CO(n379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i2 .I0_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i5  (.I0(\u_rgb2dvi/enc_0/acc[4] ), .I1(n5422), 
            .CI(n382), .O(n380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i4  (.I0(\u_rgb2dvi/enc_0/acc[3] ), .I1(n5425), 
            .CI(n384), .O(n381), .CO(n382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i3  (.I0(\u_rgb2dvi/enc_0/acc[2] ), .I1(n5428), 
            .CI(n386), .O(n383), .CO(n384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i2  (.I0(\u_rgb2dvi/enc_0/acc[1] ), .I1(n5431), 
            .CI(n3204), .O(n385), .CO(n386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_75/i5  (.I0(n366), .I1(1'b0), .CI(n353), 
            .O(n387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_0/add_75/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_75/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_75/i3  (.I0(n369), .I1(1'b0), .CI(n3048), 
            .O(n388), .CO(n389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_0/add_75/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_75/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i12  (.I0(\u_lcd_driver/vcnt[11] ), .I1(1'b0), 
            .CI(n392), .O(n390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i12 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i11  (.I0(\u_lcd_driver/vcnt[10] ), .I1(1'b0), 
            .CI(n394), .O(n391), .CO(n392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i11 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i10  (.I0(\u_lcd_driver/vcnt[9] ), .I1(1'b0), 
            .CI(n396), .O(n393), .CO(n394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i10 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i9  (.I0(\u_lcd_driver/vcnt[8] ), .I1(1'b0), 
            .CI(n398), .O(n395), .CO(n396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i9 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i8  (.I0(\u_lcd_driver/vcnt[7] ), .I1(1'b0), 
            .CI(n400), .O(n397), .CO(n398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i8 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i7  (.I0(\u_lcd_driver/vcnt[6] ), .I1(1'b0), 
            .CI(n402), .O(n399), .CO(n400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i7 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i6  (.I0(\u_lcd_driver/vcnt[5] ), .I1(1'b0), 
            .CI(n404), .O(n401), .CO(n402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i6 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i5  (.I0(\u_lcd_driver/vcnt[4] ), .I1(1'b0), 
            .CI(n406), .O(n403), .CO(n404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i5 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i4  (.I0(\u_lcd_driver/vcnt[3] ), .I1(1'b0), 
            .CI(n408), .O(n405), .CO(n406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i4 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i3  (.I0(\u_lcd_driver/vcnt[2] ), .I1(1'b0), 
            .CI(n3040), .O(n407), .CO(n408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i3 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i12  (.I0(\u_lcd_driver/hcnt[11] ), .I1(1'b0), 
            .CI(n411), .O(n409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i12 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i11  (.I0(\u_lcd_driver/hcnt[10] ), .I1(1'b0), 
            .CI(n413), .O(n410), .CO(n411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i11 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i10  (.I0(\u_lcd_driver/hcnt[9] ), .I1(1'b0), 
            .CI(n415), .O(n412), .CO(n413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i10 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i9  (.I0(\u_lcd_driver/hcnt[8] ), .I1(1'b0), 
            .CI(n417), .O(n414), .CO(n415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i9 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i8  (.I0(\u_lcd_driver/hcnt[7] ), .I1(1'b0), 
            .CI(n419), .O(n416), .CO(n417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i8 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i7  (.I0(\u_lcd_driver/hcnt[6] ), .I1(1'b0), 
            .CI(n421), .O(n418), .CO(n419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i7 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i6  (.I0(\u_lcd_driver/hcnt[5] ), .I1(1'b0), 
            .CI(n423), .O(n420), .CO(n421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i6 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i5  (.I0(\u_lcd_driver/hcnt[4] ), .I1(1'b0), 
            .CI(n425), .O(n422), .CO(n423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i5 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i4  (.I0(\u_lcd_driver/hcnt[3] ), .I1(1'b0), 
            .CI(n427), .O(n424), .CO(n425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i4 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i3  (.I0(\u_lcd_driver/hcnt[2] ), .I1(1'b0), 
            .CI(n2544), .O(n426), .CO(n427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i3 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i8  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] ), 
            .CI(n430), .O(n428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i7  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] ), 
            .CI(n432), .O(n429), .CO(n430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i6  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] ), 
            .CI(n434), .O(n431), .CO(n432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i5  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .CI(n436), .O(n433), .CO(n434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i4  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .CI(n438), .O(n435), .CO(n436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i3  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .CI(n440), .O(n437), .CO(n438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i2  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .CI(n2527), .O(n439), .CO(n440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i2  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[1] ), 
            .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[0] ), .CI(1'b0), .O(n445), 
            .CO(n446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i2 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i13  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] ), 
            .I1(1'b0), .CI(n455), .O(n453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i12  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] ), 
            .I1(1'b0), .CI(n462), .O(n454), .CO(n455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i11  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), 
            .I1(1'b0), .CI(n532), .O(n461), .CO(n462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i10  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), 
            .I1(1'b0), .CI(n542), .O(n531), .CO(n532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i9  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
            .I1(1'b0), .CI(n544), .O(n541), .CO(n542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i8  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I1(1'b0), .CI(n546), .O(n543), .CO(n544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i7  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I1(1'b0), .CI(n548), .O(n545), .CO(n546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i6  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I1(1'b0), .CI(n550), .O(n547), .CO(n548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i5  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I1(1'b0), .CI(n552), .O(n549), .CO(n550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i4  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] ), 
            .I1(1'b0), .CI(n554), .O(n551), .CO(n552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i3  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] ), 
            .I1(1'b0), .CI(n2524), .O(n553), .CO(n554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i9  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I1(1'b0), .CI(n557), .O(n555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i8  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(1'b0), .CI(n559), .O(n556), .CO(n557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i7  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(1'b0), .CI(n561), .O(n558), .CO(n559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i6  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(1'b0), .CI(n563), .O(n560), .CO(n561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i5  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(1'b0), .CI(n565), .O(n562), .CO(n563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i4  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(1'b0), .CI(n2520), .O(n564), .CO(n565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] ), 
            .I1(n5623), .CI(n568), .O(n566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] ), 
            .I1(n5626), .CI(n600), .O(n567), .CO(n568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i2  (.I0(\u_sensor_frame_count/delay_cnt[1] ), 
            .I1(\u_sensor_frame_count/delay_cnt[0] ), .CI(1'b0), .O(n575), 
            .CO(n576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i2 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] ), 
            .I1(n5660), .CI(n636), .CO(n600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i2  (.I0(\u_sensor_frame_count/cmos_fps_cnt[1] ), 
            .I1(\u_sensor_frame_count/cmos_fps_cnt[0] ), .CI(1'b0), .O(n601), 
            .CO(n602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i2 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .I1(n5723), .CI(n646), .CO(n636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i4  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .I1(n5734), .CI(n648), .CO(n646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i3  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .I1(n5737), .CI(n650), .CO(n648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i2  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I1(n5740), .CI(n2374), .CO(n650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14  (.I0(1'b0), 
            .I1(1'b1), .CI(n653), .O(n651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .CI(n655), .O(n652), .CO(n653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), .CI(n657), 
            .O(n654), .CO(n655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), .CI(n659), 
            .O(n656), .CO(n657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), .CI(n661), 
            .O(n658), .CO(n659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), .CI(n663), 
            .O(n660), .CO(n661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), .CI(n665), 
            .O(n662), .CO(n663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), .CI(n667), 
            .O(n664), .CO(n665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), .CI(n2356), 
            .O(n666), .CO(n667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I1(1'b0), .CI(n670), .O(n668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I1(1'b0), .CI(n672), .O(n669), .CO(n670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I1(1'b0), .CI(n674), .O(n671), .CO(n672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I1(1'b0), .CI(n676), .O(n673), .CO(n674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I1(1'b0), .CI(n678), .O(n675), .CO(n676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), 
            .I1(1'b0), .CI(n680), .O(n677), .CO(n678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), 
            .I1(1'b0), .CI(n2351), .O(n679), .CO(n680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
            .I1(1'b0), .CI(n697), .O(n693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/waddr[0] ), .CI(1'b0), .O(n694), 
            .CO(n695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), 
            .I1(1'b0), .CI(n718), .O(n696), .CO(n697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[2] ), 
            .I1(1'b0), .CI(n695), .O(n713), .CO(n714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), 
            .I1(1'b0), .CI(n723), .O(n717), .CO(n718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[0] ), .CI(1'b0), .O(n719), 
            .CO(n720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), 
            .I1(1'b0), .CI(n727), .O(n722), .CO(n723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1  (.I0(n5807), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[0] ), .CI(n10592), .O(n724), 
            .CO(n725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), 
            .I1(1'b0), .CI(n748), .O(n726), .CO(n727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i2  (.I0(\u_scaler_gray/vs_cnt[1] ), .I1(\u_scaler_gray/vs_cnt[0] ), 
            .CI(1'b0), .O(n745), .CO(n746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(1'b0), .CI(n750), .O(n747), .CO(n748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(1'b0), .CI(n752), .O(n749), .CO(n750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(1'b0), .CI(n754), .O(n751), .CO(n752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(1'b0), .CI(n756), .O(n753), .CO(n754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(1'b0), .CI(n2341), .O(n755), .CO(n756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i14  (.I0(\u_axi4_ctrl/araddr[23] ), .I1(1'b0), 
            .CI(n779), .O(n777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i14 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i13  (.I0(\u_axi4_ctrl/araddr[22] ), .I1(1'b0), 
            .CI(n781), .O(n778), .CO(n779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i12  (.I0(\u_axi4_ctrl/araddr[21] ), .I1(1'b0), 
            .CI(n783), .O(n780), .CO(n781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i11  (.I0(\u_axi4_ctrl/araddr[20] ), .I1(1'b0), 
            .CI(n785), .O(n782), .CO(n783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i10  (.I0(\u_axi4_ctrl/araddr[19] ), .I1(1'b0), 
            .CI(n787), .O(n784), .CO(n785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i9  (.I0(\u_axi4_ctrl/araddr[18] ), .I1(1'b0), 
            .CI(n789), .O(n786), .CO(n787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i8  (.I0(\u_axi4_ctrl/araddr[17] ), .I1(1'b0), 
            .CI(n791), .O(n788), .CO(n789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i7  (.I0(\u_axi4_ctrl/araddr[16] ), .I1(1'b0), 
            .CI(n793), .O(n790), .CO(n791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i6  (.I0(\u_axi4_ctrl/araddr[15] ), .I1(1'b0), 
            .CI(n795), .O(n792), .CO(n793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i5  (.I0(\u_axi4_ctrl/araddr[14] ), .I1(1'b0), 
            .CI(n797), .O(n794), .CO(n795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i4  (.I0(\u_axi4_ctrl/araddr[13] ), .I1(1'b0), 
            .CI(n799), .O(n796), .CO(n797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i3  (.I0(\u_axi4_ctrl/araddr[12] ), .I1(1'b0), 
            .CI(n2122), .O(n798), .CO(n799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i14  (.I0(\u_axi4_ctrl/awaddr[23] ), .I1(1'b0), 
            .CI(n802), .O(n800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i14 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i13  (.I0(\u_axi4_ctrl/awaddr[22] ), .I1(1'b0), 
            .CI(n804), .O(n801), .CO(n802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i12  (.I0(\u_axi4_ctrl/awaddr[21] ), .I1(1'b0), 
            .CI(n806), .O(n803), .CO(n804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i11  (.I0(\u_axi4_ctrl/awaddr[20] ), .I1(1'b0), 
            .CI(n808), .O(n805), .CO(n806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i10  (.I0(\u_axi4_ctrl/awaddr[19] ), .I1(1'b0), 
            .CI(n810), .O(n807), .CO(n808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i9  (.I0(\u_axi4_ctrl/awaddr[18] ), .I1(1'b0), 
            .CI(n812), .O(n809), .CO(n810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i8  (.I0(\u_axi4_ctrl/awaddr[17] ), .I1(1'b0), 
            .CI(n915), .O(n811), .CO(n812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i2  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0] ), .CI(1'b0), 
            .O(n910), .CO(n911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i7  (.I0(\u_axi4_ctrl/awaddr[16] ), .I1(1'b0), 
            .CI(n919), .O(n914), .CO(n915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i2  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] ), .CI(1'b0), 
            .O(n916), .CO(n917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i6  (.I0(\u_axi4_ctrl/awaddr[15] ), .I1(1'b0), 
            .CI(n922), .O(n918), .CO(n919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i5  (.I0(\u_axi4_ctrl/awaddr[14] ), .I1(1'b0), 
            .CI(n926), .O(n921), .CO(n922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i2  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_addra[0] ), .CI(1'b0), 
            .O(n923), .CO(n924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i4  (.I0(\u_axi4_ctrl/awaddr[13] ), .I1(1'b0), 
            .CI(n929), .O(n925), .CO(n926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i3  (.I0(\u_axi4_ctrl/awaddr[12] ), .I1(1'b0), 
            .CI(n1925), .O(n928), .CO(n929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i2  (.I0(\u_scaler_gray/destx[1] ), 
            .I1(\u_scaler_gray/destx[0] ), .CI(1'b0), .O(n930), .CO(n931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21] ), 
            .I1(1'b0), .CI(n935), .O(n933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20] ), 
            .I1(1'b0), .CI(n937), .O(n934), .CO(n935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19] ), 
            .I1(1'b0), .CI(n939), .O(n936), .CO(n937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18] ), 
            .I1(1'b0), .CI(n943), .O(n938), .CO(n939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17] ), 
            .I1(1'b0), .CI(n945), .O(n942), .CO(n943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16] ), 
            .I1(1'b0), .CI(n949), .O(n944), .CO(n945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i2  (.I0(\u_scaler_gray/desty[1] ), 
            .I1(\u_scaler_gray/desty[0] ), .CI(1'b0), .O(n946), .CO(n947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15] ), 
            .I1(1'b0), .CI(n952), .O(n948), .CO(n949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14] ), 
            .I1(1'b0), .CI(n1923), .O(n951), .CO(n952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20] ), 
            .CI(n957), .O(n954), .CO(n10593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19] ), 
            .CI(n959), .O(n956), .CO(n957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18] ), 
            .CI(n961), .O(n958), .CO(n959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17] ), 
            .CI(n963), .O(n960), .CO(n961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16] ), 
            .CI(n967), .O(n962), .CO(n963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15] ), 
            .CI(n974), .O(n966), .CO(n967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14] ), 
            .CI(n976), .O(n973), .CO(n974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13] ), 
            .CI(n1011), .O(n975), .CO(n976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12] ), 
            .CI(n1013), .O(n1010), .CO(n1011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11] ), 
            .CI(n1014), .O(n1012), .CO(n1013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10] ), 
            .CI(n1015), .CO(n1014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9] ), 
            .CI(n1016), .CO(n1015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8] ), 
            .CI(n1017), .CO(n1016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7] ), 
            .CI(n1018), .CO(n1017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6] ), 
            .CI(n1019), .CO(n1018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5] ), 
            .CI(n1020), .CO(n1019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4] ), 
            .CI(n1021), .CO(n1020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3] ), 
            .CI(n1022), .CO(n1021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2] ), 
            .CI(n1023), .CO(n1022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1] ), 
            .CI(n1920), .CO(n1023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[19] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[19] ), 
            .CI(n1027), .O(n1024), .CO(n10594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[18] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[18] ), 
            .CI(n1029), .O(n1026), .CO(n1027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[17] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[17] ), 
            .CI(n1031), .O(n1028), .CO(n1029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[16] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[16] ), 
            .CI(n1033), .O(n1030), .CO(n1031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[15] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[15] ), 
            .CI(n1035), .O(n1032), .CO(n1033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[14] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[14] ), 
            .CI(n1037), .O(n1034), .CO(n1035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[13] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[13] ), 
            .CI(n1039), .O(n1036), .CO(n1037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[12] ), 
            .CI(n1041), .O(n1038), .CO(n1039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[11] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[11] ), 
            .CI(n1043), .O(n1040), .CO(n1041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[10] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[10] ), 
            .CI(n1045), .O(n1042), .CO(n1043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[9] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[9] ), 
            .CI(n1047), .O(n1044), .CO(n1045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[8] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[8] ), 
            .CI(n1064), .O(n1046), .CO(n1047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[7] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[7] ), 
            .CI(n1066), .O(n1063), .CO(n1064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[6] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[6] ), 
            .CI(n1068), .O(n1065), .CO(n1066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[5] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[5] ), 
            .CI(n1070), .O(n1067), .CO(n1068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[4] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[4] ), 
            .CI(n1072), .O(n1069), .CO(n1070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[3] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[3] ), 
            .CI(n1074), .O(n1071), .CO(n1072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[2] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[2] ), 
            .CI(n1076), .O(n1073), .CO(n1074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[1] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[1] ), 
            .CI(n1919), .O(n1075), .CO(n1076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[19] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[19] ), 
            .CI(n1080), .O(n1077), .CO(n10595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[18] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[18] ), 
            .CI(n1082), .O(n1079), .CO(n1080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[17] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[17] ), 
            .CI(n1084), .O(n1081), .CO(n1082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[16] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[16] ), 
            .CI(n1086), .O(n1083), .CO(n1084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[15] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[15] ), 
            .CI(n1088), .O(n1085), .CO(n1086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[14] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[14] ), 
            .CI(n1090), .O(n1087), .CO(n1088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[13] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[13] ), 
            .CI(n1092), .O(n1089), .CO(n1090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[12] ), 
            .CI(n1094), .O(n1091), .CO(n1092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[11] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[11] ), 
            .CI(n1096), .O(n1093), .CO(n1094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[10] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[10] ), 
            .CI(n1098), .O(n1095), .CO(n1096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[9] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[9] ), 
            .CI(n1100), .O(n1097), .CO(n1098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[8] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[8] ), 
            .CI(n1102), .O(n1099), .CO(n1100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[7] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[7] ), 
            .CI(n1104), .O(n1101), .CO(n1102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[6] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[6] ), 
            .CI(n1106), .O(n1103), .CO(n1104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[5] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[5] ), 
            .CI(n1108), .O(n1105), .CO(n1106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[4] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[4] ), 
            .CI(n1110), .O(n1107), .CO(n1108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[3] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[3] ), 
            .CI(n1114), .O(n1109), .CO(n1110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[2] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[2] ), 
            .CI(n1116), .O(n1113), .CO(n1114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[1] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[1] ), 
            .CI(n1754), .O(n1115), .CO(n1116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[23] ), 
            .I1(1'b0), .CI(n1135), .O(n1133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[22] ), 
            .I1(1'b0), .CI(n1137), .O(n1134), .CO(n1135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[21] ), 
            .I1(1'b0), .CI(n1139), .O(n1136), .CO(n1137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[20] ), 
            .I1(1'b0), .CI(n1141), .O(n1138), .CO(n1139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[19] ), 
            .I1(1'b0), .CI(n1143), .O(n1140), .CO(n1141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[18] ), 
            .I1(1'b0), .CI(n1145), .O(n1142), .CO(n1143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[17] ), 
            .I1(1'b0), .CI(n1147), .O(n1144), .CO(n1145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[16] ), 
            .I1(1'b0), .CI(n1149), .O(n1146), .CO(n1147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[15] ), 
            .I1(1'b0), .CI(n1151), .O(n1148), .CO(n1149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[14] ), 
            .I1(1'b0), .CI(n1153), .O(n1150), .CO(n1151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[13] ), 
            .I1(1'b0), .CI(n1736), .O(n1152), .CO(n1153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[23] ), 
            .I1(1'b0), .CI(n1156), .O(n1154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[22] ), 
            .I1(1'b0), .CI(n1158), .O(n1155), .CO(n1156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[21] ), 
            .I1(1'b0), .CI(n1160), .O(n1157), .CO(n1158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[20] ), 
            .I1(1'b0), .CI(n1162), .O(n1159), .CO(n1160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[19] ), 
            .I1(1'b0), .CI(n1164), .O(n1161), .CO(n1162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[18] ), 
            .I1(1'b0), .CI(n1166), .O(n1163), .CO(n1164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[17] ), 
            .I1(1'b0), .CI(n1168), .O(n1165), .CO(n1166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[16] ), 
            .I1(1'b0), .CI(n1170), .O(n1167), .CO(n1168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[15] ), 
            .I1(1'b0), .CI(n1172), .O(n1169), .CO(n1170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[14] ), 
            .I1(1'b0), .CI(n1174), .O(n1171), .CO(n1172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[13] ), 
            .I1(1'b0), .CI(n1734), .O(n1173), .CO(n1174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[23] ), 
            .I1(1'b0), .CI(n1177), .O(n1175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[22] ), 
            .I1(1'b0), .CI(n1179), .O(n1176), .CO(n1177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[21] ), 
            .I1(1'b0), .CI(n1181), .O(n1178), .CO(n1179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[20] ), 
            .I1(1'b0), .CI(n1183), .O(n1180), .CO(n1181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[19] ), 
            .I1(1'b0), .CI(n1200), .O(n1182), .CO(n1183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[18] ), 
            .I1(1'b0), .CI(n1202), .O(n1199), .CO(n1200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[17] ), 
            .I1(1'b0), .CI(n1204), .O(n1201), .CO(n1202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[16] ), 
            .I1(1'b0), .CI(n1206), .O(n1203), .CO(n1204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[15] ), 
            .I1(1'b0), .CI(n1208), .O(n1205), .CO(n1206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[14] ), 
            .I1(1'b0), .CI(n1210), .O(n1207), .CO(n1208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[13] ), 
            .I1(1'b0), .CI(n1732), .O(n1209), .CO(n1210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[23] ), 
            .I1(1'b0), .CI(n1213), .O(n1211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[22] ), 
            .I1(1'b0), .CI(n1215), .O(n1212), .CO(n1213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[21] ), 
            .I1(1'b0), .CI(n1217), .O(n1214), .CO(n1215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[20] ), 
            .I1(1'b0), .CI(n1219), .O(n1216), .CO(n1217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[19] ), 
            .I1(1'b0), .CI(n1221), .O(n1218), .CO(n1219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[18] ), 
            .I1(1'b0), .CI(n1223), .O(n1220), .CO(n1221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[17] ), 
            .I1(1'b0), .CI(n1225), .O(n1222), .CO(n1223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[16] ), 
            .I1(1'b0), .CI(n1227), .O(n1224), .CO(n1225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[15] ), 
            .I1(1'b0), .CI(n1229), .O(n1226), .CO(n1227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[14] ), 
            .I1(1'b0), .CI(n1231), .O(n1228), .CO(n1229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[13] ), 
            .I1(1'b0), .CI(n1689), .O(n1230), .CO(n1231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i28  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27] ), 
            .I1(1'b1), .CI(n1234), .O(n1232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i27  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26] ), 
            .I1(1'b1), .CI(n1236), .O(n1233), .CO(n1234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i26  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25] ), 
            .I1(1'b1), .CI(n1238), .O(n1235), .CO(n1236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i25  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24] ), 
            .I1(1'b1), .CI(n1240), .O(n1237), .CO(n1238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i24  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23] ), 
            .I1(1'b1), .CI(n1242), .O(n1239), .CO(n1240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i23  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22] ), 
            .I1(1'b1), .CI(n1244), .O(n1241), .CO(n1242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i22  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21] ), 
            .I1(1'b1), .CI(n1246), .O(n1243), .CO(n1244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i21  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20] ), 
            .I1(1'b1), .CI(n1248), .O(n1245), .CO(n1246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19] ), 
            .I1(1'b1), .CI(n1250), .O(n1247), .CO(n1248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18] ), 
            .I1(1'b1), .CI(n1252), .O(n1249), .CO(n1250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17] ), 
            .I1(1'b1), .CI(n1254), .O(n1251), .CO(n1252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16] ), 
            .I1(1'b1), .CI(n1256), .O(n1253), .CO(n1254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15] ), 
            .I1(1'b1), .CI(n1258), .O(n1255), .CO(n1256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14] ), 
            .I1(1'b1), .CI(n1260), .O(n1257), .CO(n1258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13] ), 
            .I1(1'b1), .CI(n1262), .O(n1259), .CO(n1260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12] ), 
            .I1(1'b1), .CI(n1687), .O(n1261), .CO(n1262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i28  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27] ), 
            .CI(n1265), .O(n1263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i27  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26] ), 
            .CI(n1267), .O(n1264), .CO(n1265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i26  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25] ), 
            .CI(n1273), .O(n1266), .CO(n1267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i25  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24] ), 
            .CI(n1275), .O(n1272), .CO(n1273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i24  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23] ), 
            .CI(n1277), .O(n1274), .CO(n1275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i23  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22] ), 
            .CI(n1279), .O(n1276), .CO(n1277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i22  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21] ), 
            .CI(n1281), .O(n1278), .CO(n1279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i21  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20] ), 
            .CI(n1283), .O(n1280), .CO(n1281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i20  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19] ), 
            .CI(n1285), .O(n1282), .CO(n1283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i19  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18] ), 
            .CI(n1287), .O(n1284), .CO(n1285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i18  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17] ), 
            .CI(n1289), .O(n1286), .CO(n1287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i17  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16] ), 
            .CI(n1291), .O(n1288), .CO(n1289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i16  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15] ), 
            .CI(n1293), .O(n1290), .CO(n1291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i15  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14] ), 
            .CI(n1295), .O(n1292), .CO(n1293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i14  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13] ), 
            .CI(n1297), .O(n1294), .CO(n1295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i13  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12] ), 
            .CI(n1299), .O(n1296), .CO(n1297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i12  (.I0(1'b1), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11] ), 
            .CI(n1301), .O(n1298), .CO(n1299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i11  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10] ), 
            .CI(n1303), .O(n1300), .CO(n1301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i10  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9] ), 
            .CI(n1305), .O(n1302), .CO(n1303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i9  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8] ), 
            .CI(n1307), .O(n1304), .CO(n1305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i8  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7] ), 
            .CI(n1309), .O(n1306), .CO(n1307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i7  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6] ), 
            .CI(n1311), .O(n1308), .CO(n1309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i6  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5] ), 
            .CI(n1313), .O(n1310), .CO(n1311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i5  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4] ), 
            .CI(n1315), .O(n1312), .CO(n1313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i4  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3] ), 
            .CI(n1317), .O(n1314), .CO(n1315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i3  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2] ), 
            .CI(n1319), .O(n1316), .CO(n1317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i2  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1] ), 
            .CI(n1657), .O(n1318), .CO(n1319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i28  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27] ), 
            .I1(1'b1), .CI(n1322), .O(n1320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i27  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26] ), 
            .I1(1'b1), .CI(n1324), .O(n1321), .CO(n1322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i26  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25] ), 
            .I1(1'b1), .CI(n1326), .O(n1323), .CO(n1324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i25  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24] ), 
            .I1(1'b1), .CI(n1328), .O(n1325), .CO(n1326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i24  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23] ), 
            .I1(1'b1), .CI(n1330), .O(n1327), .CO(n1328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i23  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22] ), 
            .I1(1'b1), .CI(n1332), .O(n1329), .CO(n1330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i22  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21] ), 
            .I1(1'b1), .CI(n1334), .O(n1331), .CO(n1332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i21  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20] ), 
            .I1(1'b1), .CI(n1336), .O(n1333), .CO(n1334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19] ), 
            .I1(1'b1), .CI(n1338), .O(n1335), .CO(n1336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18] ), 
            .I1(1'b1), .CI(n1340), .O(n1337), .CO(n1338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17] ), 
            .I1(1'b1), .CI(n1364), .O(n1339), .CO(n1340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16] ), 
            .I1(1'b1), .CI(n1366), .O(n1363), .CO(n1364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15] ), 
            .I1(1'b1), .CI(n1368), .O(n1365), .CO(n1366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14] ), 
            .I1(1'b1), .CI(n1370), .O(n1367), .CO(n1368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13] ), 
            .I1(1'b1), .CI(n1372), .O(n1369), .CO(n1370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12] ), 
            .I1(1'b1), .CI(n1655), .O(n1371), .CO(n1372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i28  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27] ), 
            .CI(n1412), .O(n1410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i27  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26] ), 
            .CI(n1414), .O(n1411), .CO(n1412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i26  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25] ), 
            .CI(n1416), .O(n1413), .CO(n1414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i25  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24] ), 
            .CI(n1418), .O(n1415), .CO(n1416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i24  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23] ), 
            .CI(n1420), .O(n1417), .CO(n1418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i23  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22] ), 
            .CI(n1464), .O(n1419), .CO(n1420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i22  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21] ), 
            .CI(n1466), .O(n1463), .CO(n1464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i21  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20] ), 
            .CI(n1468), .O(n1465), .CO(n1466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i20  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19] ), 
            .CI(n1470), .O(n1467), .CO(n1468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i19  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18] ), 
            .CI(n1472), .O(n1469), .CO(n1470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i18  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17] ), 
            .CI(n1474), .O(n1471), .CO(n1472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i17  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16] ), 
            .CI(n1476), .O(n1473), .CO(n1474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i16  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15] ), 
            .CI(n1478), .O(n1475), .CO(n1476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i15  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14] ), 
            .CI(n1480), .O(n1477), .CO(n1478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i14  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13] ), 
            .CI(n1482), .O(n1479), .CO(n1480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i13  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12] ), 
            .CI(n1484), .O(n1481), .CO(n1482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i12  (.I0(1'b1), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11] ), 
            .CI(n1486), .O(n1483), .CO(n1484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i11  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10] ), 
            .CI(n1488), .O(n1485), .CO(n1486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10  (.I0(1'b0), 
            .I1(DdrCtrl_ALEN_0[0]), .CI(n10596), .O(n1487), .CO(n1488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \add_344/i28  (.I0(1'b0), .I1(\u_scaler_gray/destx[15] ), .CI(n1491), 
            .O(n1489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i28 .I0_POLARITY = 1'b1;
    defparam \add_344/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i27  (.I0(1'b0), .I1(\u_scaler_gray/destx[14] ), .CI(n1493), 
            .O(n1490), .CO(n1491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i27 .I0_POLARITY = 1'b1;
    defparam \add_344/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i26  (.I0(\u_scaler_gray/destx[15] ), .I1(\u_scaler_gray/destx[13] ), 
            .CI(n1495), .O(n1492), .CO(n1493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i26 .I0_POLARITY = 1'b1;
    defparam \add_344/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i25  (.I0(\u_scaler_gray/destx[14] ), .I1(\u_scaler_gray/destx[12] ), 
            .CI(n1497), .O(n1494), .CO(n1495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i25 .I0_POLARITY = 1'b1;
    defparam \add_344/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i24  (.I0(\u_scaler_gray/destx[13] ), .I1(\u_scaler_gray/destx[11] ), 
            .CI(n1499), .O(n1496), .CO(n1497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i24 .I0_POLARITY = 1'b1;
    defparam \add_344/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i23  (.I0(\u_scaler_gray/destx[12] ), .I1(\u_scaler_gray/destx[10] ), 
            .CI(n1501), .O(n1498), .CO(n1499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i23 .I0_POLARITY = 1'b1;
    defparam \add_344/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i22  (.I0(\u_scaler_gray/destx[11] ), .I1(\u_scaler_gray/destx[9] ), 
            .CI(n1503), .O(n1500), .CO(n1501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i22 .I0_POLARITY = 1'b1;
    defparam \add_344/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i21  (.I0(\u_scaler_gray/destx[10] ), .I1(\u_scaler_gray/destx[8] ), 
            .CI(n1505), .O(n1502), .CO(n1503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i21 .I0_POLARITY = 1'b1;
    defparam \add_344/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i20  (.I0(\u_scaler_gray/destx[9] ), .I1(\u_scaler_gray/destx[7] ), 
            .CI(n1507), .O(n1504), .CO(n1505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i20 .I0_POLARITY = 1'b1;
    defparam \add_344/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i19  (.I0(\u_scaler_gray/destx[8] ), .I1(\u_scaler_gray/destx[6] ), 
            .CI(n1509), .O(n1506), .CO(n1507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i19 .I0_POLARITY = 1'b1;
    defparam \add_344/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i18  (.I0(\u_scaler_gray/destx[7] ), .I1(\u_scaler_gray/destx[5] ), 
            .CI(n1511), .O(n1508), .CO(n1509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i18 .I0_POLARITY = 1'b1;
    defparam \add_344/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i17  (.I0(\u_scaler_gray/destx[6] ), .I1(\u_scaler_gray/destx[4] ), 
            .CI(n1513), .O(n1510), .CO(n1511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i17 .I0_POLARITY = 1'b1;
    defparam \add_344/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i16  (.I0(\u_scaler_gray/destx[5] ), .I1(\u_scaler_gray/destx[3] ), 
            .CI(n1515), .O(n1512), .CO(n1513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i16 .I0_POLARITY = 1'b1;
    defparam \add_344/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i15  (.I0(\u_scaler_gray/destx[4] ), .I1(\u_scaler_gray/destx[2] ), 
            .CI(n1517), .O(n1514), .CO(n1515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i15 .I0_POLARITY = 1'b1;
    defparam \add_344/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i14  (.I0(\u_scaler_gray/destx[3] ), .I1(\u_scaler_gray/destx[1] ), 
            .CI(n1538), .O(n1516), .CO(n1517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i14 .I0_POLARITY = 1'b1;
    defparam \add_344/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[1] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[0] ), 
            .CI(1'b0), .O(n1535), .CO(n1536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_344/i13  (.I0(\u_scaler_gray/destx[2] ), .I1(\u_scaler_gray/destx[0] ), 
            .CI(1'b0), .O(n1537), .CO(n1538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_344/i13 .I0_POLARITY = 1'b1;
    defparam \add_344/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11] ), 
            .I1(1'b0), .CI(n10597), .O(n1654), .CO(n1655)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0] ), 
            .CI(n10598), .O(n1656), .CO(n1657)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i28  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[27] ), 
            .I1(1'b0), .CI(n1691), .O(n1685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11] ), 
            .I1(1'b0), .CI(n10599), .O(n1686), .CO(n1687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[11] ), 
            .CI(1'b0), .O(n1688), .CO(n1689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i27  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[26] ), 
            .I1(1'b0), .CI(n1693), .O(n1690), .CO(n1691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i26  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[25] ), 
            .I1(1'b0), .CI(n1695), .O(n1692), .CO(n1693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i25  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[24] ), 
            .I1(1'b0), .CI(n1697), .O(n1694), .CO(n1695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i24  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[23] ), 
            .I1(1'b0), .CI(n1699), .O(n1696), .CO(n1697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i23  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[22] ), 
            .I1(1'b0), .CI(n1701), .O(n1698), .CO(n1699)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i22  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[21] ), 
            .I1(1'b0), .CI(n1703), .O(n1700), .CO(n1701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i21  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[20] ), 
            .I1(1'b0), .CI(n1705), .O(n1702), .CO(n1703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[19] ), 
            .I1(1'b0), .CI(n1707), .O(n1704), .CO(n1705)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[18] ), 
            .I1(1'b0), .CI(n1741), .O(n1706), .CO(n1707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[11] ), 
            .CI(1'b0), .O(n1731), .CO(n1732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[11] ), 
            .CI(1'b0), .O(n1733), .CO(n1734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[11] ), 
            .CI(1'b0), .O(n1735), .CO(n1736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[17] ), 
            .I1(1'b0), .CI(n1784), .O(n1740), .CO(n1741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[0] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[0] ), 
            .CI(1'b0), .O(n1753), .CO(n1754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[16] ), 
            .I1(1'b0), .CI(n2055), .O(n1783), .CO(n1784)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[0] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[0] ), 
            .CI(1'b0), .O(n1918), .CO(n1919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0] ), 
            .CI(1'b0), .CO(n1920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12] ), 
            .CI(1'b0), .O(n1922), .CO(n1923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i2  (.I0(\u_axi4_ctrl/awaddr[11] ), .I1(\u_axi4_ctrl/awaddr[10] ), 
            .CI(1'b0), .O(n1924), .CO(n1925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[15] ), 
            .I1(1'b0), .CI(n2057), .O(n2054), .CO(n2055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[14] ), 
            .I1(1'b0), .CI(n2059), .O(n2056), .CO(n2057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[13] ), 
            .I1(1'b0), .CI(n2061), .O(n2058), .CO(n2059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[12] ), 
            .I1(1'b0), .CI(n2063), .O(n2060), .CO(n2061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[11] ), 
            .I1(1'b1), .CI(n2065), .O(n2062), .CO(n2063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[10] ), 
            .I1(1'b0), .CI(n2067), .O(n2064), .CO(n2065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[9] ), 
            .I1(1'b0), .CI(n2092), .O(n2066), .CO(n2067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[8] ), 
            .I1(1'b1), .CI(n2094), .O(n2091), .CO(n2092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[7] ), 
            .I1(1'b1), .CI(n2097), .O(n2093), .CO(n2094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[6] ), 
            .I1(1'b0), .CI(n2099), .O(n2096), .CO(n2097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[5] ), 
            .I1(1'b0), .CI(n2103), .O(n2098), .CO(n2099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[4] ), 
            .I1(1'b1), .CI(n2106), .O(n2102), .CO(n2103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[3] ), 
            .I1(1'b1), .CI(n2108), .O(n2105), .CO(n2106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[2] ), 
            .I1(1'b0), .CI(n1536), .O(n2107), .CO(n2108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i28  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27] ), 
            .I1(1'b0), .CI(n2113), .O(n2110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i27  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26] ), 
            .I1(1'b0), .CI(n2116), .O(n2112), .CO(n2113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i26  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25] ), 
            .I1(1'b0), .CI(n2118), .O(n2115), .CO(n2116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i25  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24] ), 
            .I1(1'b0), .CI(n2120), .O(n2117), .CO(n2118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i24  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23] ), 
            .I1(1'b0), .CI(n2124), .O(n2119), .CO(n2120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i2  (.I0(\u_axi4_ctrl/araddr[11] ), .I1(\u_axi4_ctrl/araddr[10] ), 
            .CI(1'b0), .O(n2121), .CO(n2122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i23  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22] ), 
            .I1(1'b0), .CI(n2126), .O(n2123), .CO(n2124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i22  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21] ), 
            .I1(1'b0), .CI(n2130), .O(n2125), .CO(n2126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i21  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20] ), 
            .I1(1'b0), .CI(n2135), .O(n2129), .CO(n2130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19] ), 
            .I1(1'b0), .CI(n2137), .O(n2134), .CO(n2135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18] ), 
            .I1(1'b0), .CI(n2139), .O(n2136), .CO(n2137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17] ), 
            .I1(1'b0), .CI(n2141), .O(n2138), .CO(n2139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16] ), 
            .I1(1'b0), .CI(n2143), .O(n2140), .CO(n2141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15] ), 
            .I1(1'b0), .CI(n2147), .O(n2142), .CO(n2143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14] ), 
            .I1(1'b0), .CI(n2149), .O(n2146), .CO(n2147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13] ), 
            .I1(1'b0), .CI(n2151), .O(n2148), .CO(n2149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12] ), 
            .I1(1'b0), .CI(n2153), .O(n2150), .CO(n2151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11] ), 
            .I1(1'b1), .CI(1'b0), .O(n2152), .CO(n2153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i16  (.I0(\u_scaler_gray/desty[15] ), 
            .I1(1'b0), .CI(n2156), .O(n2154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i15  (.I0(\u_scaler_gray/desty[14] ), 
            .I1(1'b0), .CI(n2158), .O(n2155), .CO(n2156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i14  (.I0(\u_scaler_gray/desty[13] ), 
            .I1(1'b0), .CI(n2160), .O(n2157), .CO(n2158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i13  (.I0(\u_scaler_gray/desty[12] ), 
            .I1(1'b0), .CI(n2162), .O(n2159), .CO(n2160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i12  (.I0(\u_scaler_gray/desty[11] ), 
            .I1(1'b0), .CI(n2164), .O(n2161), .CO(n2162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i11  (.I0(\u_scaler_gray/desty[10] ), 
            .I1(1'b0), .CI(n2166), .O(n2163), .CO(n2164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i10  (.I0(\u_scaler_gray/desty[9] ), 
            .I1(1'b0), .CI(n2168), .O(n2165), .CO(n2166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i9  (.I0(\u_scaler_gray/desty[8] ), 
            .I1(1'b0), .CI(n2170), .O(n2167), .CO(n2168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i8  (.I0(\u_scaler_gray/desty[7] ), 
            .I1(1'b0), .CI(n2172), .O(n2169), .CO(n2170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i7  (.I0(\u_scaler_gray/desty[6] ), 
            .I1(1'b0), .CI(n2174), .O(n2171), .CO(n2172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i6  (.I0(\u_scaler_gray/desty[5] ), 
            .I1(1'b0), .CI(n2176), .O(n2173), .CO(n2174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i5  (.I0(\u_scaler_gray/desty[4] ), 
            .I1(1'b0), .CI(n2178), .O(n2175), .CO(n2176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i4  (.I0(\u_scaler_gray/desty[3] ), 
            .I1(1'b0), .CI(n2180), .O(n2177), .CO(n2178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i3  (.I0(\u_scaler_gray/desty[2] ), 
            .I1(1'b0), .CI(n947), .O(n2179), .CO(n2180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i16  (.I0(\u_scaler_gray/destx[15] ), 
            .I1(1'b0), .CI(n2186), .O(n2184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i15  (.I0(\u_scaler_gray/destx[14] ), 
            .I1(1'b0), .CI(n2188), .O(n2185), .CO(n2186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i14  (.I0(\u_scaler_gray/destx[13] ), 
            .I1(1'b0), .CI(n2190), .O(n2187), .CO(n2188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i13  (.I0(\u_scaler_gray/destx[12] ), 
            .I1(1'b0), .CI(n2215), .O(n2189), .CO(n2190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i12  (.I0(\u_scaler_gray/destx[11] ), 
            .I1(1'b0), .CI(n2217), .O(n2214), .CO(n2215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i11  (.I0(\u_scaler_gray/destx[10] ), 
            .I1(1'b0), .CI(n2219), .O(n2216), .CO(n2217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i10  (.I0(\u_scaler_gray/destx[9] ), 
            .I1(1'b0), .CI(n2221), .O(n2218), .CO(n2219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i9  (.I0(\u_scaler_gray/destx[8] ), 
            .I1(1'b0), .CI(n2347), .O(n2220), .CO(n2221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] ), .CI(1'b0), 
            .O(n2322), .CO(n2323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(1'b0), .CI(n2323), .O(n2340), .CO(n2341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i8  (.I0(\u_scaler_gray/destx[7] ), 
            .I1(1'b0), .CI(n2349), .O(n2346), .CO(n2347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i7  (.I0(\u_scaler_gray/destx[6] ), 
            .I1(1'b0), .CI(n2354), .O(n2348), .CO(n2349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), .CI(1'b0), 
            .O(n2350), .CO(n2351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i6  (.I0(\u_scaler_gray/destx[5] ), 
            .I1(1'b0), .CI(n2358), .O(n2353), .CO(n2354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), .CI(n10601), 
            .O(n2355), .CO(n2356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i5  (.I0(\u_scaler_gray/destx[4] ), 
            .I1(1'b0), .CI(n2377), .O(n2357), .CO(n2358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .I1(n7366), .CI(n10602), .CO(n2374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i4  (.I0(\u_scaler_gray/destx[3] ), 
            .I1(1'b0), .CI(n2379), .O(n2376), .CO(n2377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i3  (.I0(\u_scaler_gray/destx[2] ), 
            .I1(1'b0), .CI(n931), .O(n2378), .CO(n2379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i16  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[15] ), 
            .I1(1'b0), .CI(n2382), .O(n2380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i15  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[14] ), 
            .I1(1'b0), .CI(n2384), .O(n2381), .CO(n2382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i14  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[13] ), 
            .I1(1'b0), .CI(n2386), .O(n2383), .CO(n2384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i13  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[12] ), 
            .I1(1'b0), .CI(n2388), .O(n2385), .CO(n2386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i12  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[11] ), 
            .I1(1'b0), .CI(n2398), .O(n2387), .CO(n2388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i11  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[10] ), 
            .I1(1'b0), .CI(n2400), .O(n2397), .CO(n2398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i10  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[9] ), 
            .I1(1'b0), .CI(n2402), .O(n2399), .CO(n2400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i9  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[8] ), 
            .I1(1'b0), .CI(n2404), .O(n2401), .CO(n2402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i8  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[7] ), 
            .I1(1'b0), .CI(n2406), .O(n2403), .CO(n2404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i7  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[6] ), 
            .I1(1'b0), .CI(n2408), .O(n2405), .CO(n2406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i6  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[5] ), 
            .I1(1'b0), .CI(n2489), .O(n2407), .CO(n2408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i5  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[4] ), 
            .I1(1'b0), .CI(n2491), .O(n2488), .CO(n2489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i4  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[3] ), 
            .I1(1'b0), .CI(n2493), .O(n2490), .CO(n2491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i3  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[2] ), 
            .I1(1'b0), .CI(n924), .O(n2492), .CO(n2493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i16  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] ), 
            .I1(1'b0), .CI(n2496), .O(n2494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i15  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] ), 
            .I1(1'b0), .CI(n2498), .O(n2495), .CO(n2496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i14  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] ), 
            .I1(1'b0), .CI(n2500), .O(n2497), .CO(n2498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i13  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] ), 
            .I1(1'b0), .CI(n2502), .O(n2499), .CO(n2500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i12  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] ), 
            .I1(1'b0), .CI(n2504), .O(n2501), .CO(n2502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i11  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] ), 
            .I1(1'b0), .CI(n2506), .O(n2503), .CO(n2504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i10  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] ), 
            .I1(1'b0), .CI(n2529), .O(n2505), .CO(n2506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i2  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), .CI(1'b0), 
            .O(n2516), .CO(n2517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i3  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(1'b0), .CI(n2517), .O(n2519), .CO(n2520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i2  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] ), .CI(1'b0), 
            .O(n2523), .CO(n2524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .CI(n10603), .O(n2526), .CO(n2527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i9  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] ), 
            .I1(1'b0), .CI(n2534), .O(n2528), .CO(n2529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i8  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] ), 
            .I1(1'b0), .CI(n2546), .O(n2533), .CO(n2534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i2  (.I0(\u_lcd_driver/hcnt[1] ), .I1(\u_lcd_driver/hcnt[0] ), 
            .CI(1'b0), .O(n2543), .CO(n2544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i2 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i7  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] ), 
            .I1(1'b0), .CI(n2548), .O(n2545), .CO(n2546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i6  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] ), 
            .I1(1'b0), .CI(n2550), .O(n2547), .CO(n2548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i5  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] ), 
            .I1(1'b0), .CI(n2552), .O(n2549), .CO(n2550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i4  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] ), 
            .I1(1'b0), .CI(n2554), .O(n2551), .CO(n2552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i3  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] ), 
            .I1(1'b0), .CI(n917), .O(n2553), .CO(n2554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i16  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15] ), 
            .I1(1'b0), .CI(n2569), .O(n2555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i15  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14] ), 
            .I1(1'b0), .CI(n2571), .O(n2568), .CO(n2569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i14  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13] ), 
            .I1(1'b0), .CI(n2573), .O(n2570), .CO(n2571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i13  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12] ), 
            .I1(1'b0), .CI(n2575), .O(n2572), .CO(n2573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i12  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11] ), 
            .I1(1'b0), .CI(n2577), .O(n2574), .CO(n2575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i11  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10] ), 
            .I1(1'b0), .CI(n2579), .O(n2576), .CO(n2577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i10  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9] ), 
            .I1(1'b0), .CI(n2581), .O(n2578), .CO(n2579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i9  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8] ), 
            .I1(1'b0), .CI(n2583), .O(n2580), .CO(n2581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i8  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7] ), 
            .I1(1'b0), .CI(n2585), .O(n2582), .CO(n2583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i7  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6] ), 
            .I1(1'b0), .CI(n2587), .O(n2584), .CO(n2585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i6  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5] ), 
            .I1(1'b0), .CI(n2589), .O(n2586), .CO(n2587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i5  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4] ), 
            .I1(1'b0), .CI(n2591), .O(n2588), .CO(n2589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i4  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3] ), 
            .I1(1'b0), .CI(n2593), .O(n2590), .CO(n2591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i3  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2] ), 
            .I1(1'b0), .CI(n911), .O(n2592), .CO(n2593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i16  (.I0(\u_scaler_gray/vs_cnt[15] ), .I1(1'b0), 
            .CI(n2596), .O(n2594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i15  (.I0(\u_scaler_gray/vs_cnt[14] ), .I1(1'b0), 
            .CI(n2598), .O(n2595), .CO(n2596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i14  (.I0(\u_scaler_gray/vs_cnt[13] ), .I1(1'b0), 
            .CI(n2600), .O(n2597), .CO(n2598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i13  (.I0(\u_scaler_gray/vs_cnt[12] ), .I1(1'b0), 
            .CI(n2602), .O(n2599), .CO(n2600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i12  (.I0(\u_scaler_gray/vs_cnt[11] ), .I1(1'b0), 
            .CI(n2604), .O(n2601), .CO(n2602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i11  (.I0(\u_scaler_gray/vs_cnt[10] ), .I1(1'b0), 
            .CI(n2606), .O(n2603), .CO(n2604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i10  (.I0(\u_scaler_gray/vs_cnt[9] ), .I1(1'b0), 
            .CI(n2688), .O(n2605), .CO(n2606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i9  (.I0(\u_scaler_gray/vs_cnt[8] ), .I1(1'b0), 
            .CI(n2690), .O(n2687), .CO(n2688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i8  (.I0(\u_scaler_gray/vs_cnt[7] ), .I1(1'b0), 
            .CI(n2692), .O(n2689), .CO(n2690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i7  (.I0(\u_scaler_gray/vs_cnt[6] ), .I1(1'b0), 
            .CI(n2695), .O(n2691), .CO(n2692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i6  (.I0(\u_scaler_gray/vs_cnt[5] ), .I1(1'b0), 
            .CI(n2697), .O(n2694), .CO(n2695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i5  (.I0(\u_scaler_gray/vs_cnt[4] ), .I1(1'b0), 
            .CI(n2701), .O(n2696), .CO(n2697)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i4  (.I0(\u_scaler_gray/vs_cnt[3] ), .I1(1'b0), 
            .CI(n2703), .O(n2700), .CO(n2701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i3  (.I0(\u_scaler_gray/vs_cnt[2] ), .I1(1'b0), 
            .CI(n746), .O(n2702), .CO(n2703)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i15  (.I0(1'b0), 
            .I1(1'b1), .CI(n2740), .O(n2738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14  (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] ), 
            .CI(n2742), .O(n2739), .CO(n2740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13  (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_q ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), .CI(n2744), .O(n2741), 
            .CO(n2742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12  (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1_q ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[11] ), .CI(n2746), .O(n2743), 
            .CO(n2744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11  (.I0(n7832), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[10] ), .CI(n2748), .O(n2745), 
            .CO(n2746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10  (.I0(n7835), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[9] ), .CI(n2750), .O(n2747), 
            .CO(n2748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9  (.I0(n7838), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[8] ), .CI(n2752), .O(n2749), 
            .CO(n2750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8  (.I0(n7841), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[7] ), .CI(n2754), .O(n2751), 
            .CO(n2752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7  (.I0(n7844), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[6] ), .CI(n2756), .O(n2753), 
            .CO(n2754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6  (.I0(n7847), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[5] ), .CI(n2758), .O(n2755), 
            .CO(n2756)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5  (.I0(n7850), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[4] ), .CI(n2760), .O(n2757), 
            .CO(n2758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4  (.I0(n7853), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[3] ), .CI(n2762), .O(n2759), 
            .CO(n2760)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i3  (.I0(n7856), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[2] ), .CI(n2764), .O(n2761), 
            .CO(n2762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i2  (.I0(n7859), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[1] ), .CI(n725), .O(n2763), 
            .CO(n2764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i14  (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] ), 
            .I1(1'b0), .CI(n2767), .O(n2765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i14 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i13  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), 
            .I1(1'b0), .CI(n2769), .O(n2766), .CO(n2767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i13 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i12  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[11] ), 
            .I1(1'b0), .CI(n2771), .O(n2768), .CO(n2769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i12 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i11  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[10] ), 
            .I1(1'b0), .CI(n2773), .O(n2770), .CO(n2771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i11 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i10  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[9] ), 
            .I1(1'b0), .CI(n2775), .O(n2772), .CO(n2773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i10 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[8] ), 
            .I1(1'b0), .CI(n2777), .O(n2774), .CO(n2775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[7] ), 
            .I1(1'b0), .CI(n2779), .O(n2776), .CO(n2777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[6] ), 
            .I1(1'b0), .CI(n2781), .O(n2778), .CO(n2779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[5] ), 
            .I1(1'b0), .CI(n2783), .O(n2780), .CO(n2781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[4] ), 
            .I1(1'b0), .CI(n2785), .O(n2782), .CO(n2783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[3] ), 
            .I1(1'b0), .CI(n2787), .O(n2784), .CO(n2785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[2] ), 
            .I1(1'b0), .CI(n720), .O(n2786), .CO(n2787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i14  (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] ), 
            .I1(1'b0), .CI(n2804), .O(n2802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i14 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), 
            .I1(1'b0), .CI(n2806), .O(n2803), .CO(n2804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[11] ), 
            .I1(1'b0), .CI(n2808), .O(n2805), .CO(n2806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[10] ), 
            .I1(1'b0), .CI(n2810), .O(n2807), .CO(n2808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[9] ), 
            .I1(1'b0), .CI(n2812), .O(n2809), .CO(n2810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[8] ), 
            .I1(1'b0), .CI(n2814), .O(n2811), .CO(n2812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[7] ), 
            .I1(1'b0), .CI(n2816), .O(n2813), .CO(n2814)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[6] ), 
            .I1(1'b0), .CI(n2818), .O(n2815), .CO(n2816)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[5] ), 
            .I1(1'b0), .CI(n2820), .O(n2817), .CO(n2818)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[4] ), 
            .I1(1'b0), .CI(n2822), .O(n2819), .CO(n2820)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[3] ), 
            .I1(1'b0), .CI(n714), .O(n2821), .CO(n2822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i9  (.I0(\u_sensor_frame_count/cmos_fps_cnt[8] ), 
            .I1(1'b0), .CI(n2867), .O(n2865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i9 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i8  (.I0(\u_sensor_frame_count/cmos_fps_cnt[7] ), 
            .I1(1'b0), .CI(n2869), .O(n2866), .CO(n2867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i8 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i7  (.I0(\u_sensor_frame_count/cmos_fps_cnt[6] ), 
            .I1(1'b0), .CI(n2871), .O(n2868), .CO(n2869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i7 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i6  (.I0(\u_sensor_frame_count/cmos_fps_cnt[5] ), 
            .I1(1'b0), .CI(n2873), .O(n2870), .CO(n2871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i6 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i5  (.I0(\u_sensor_frame_count/cmos_fps_cnt[4] ), 
            .I1(1'b0), .CI(n2875), .O(n2872), .CO(n2873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i5 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i4  (.I0(\u_sensor_frame_count/cmos_fps_cnt[3] ), 
            .I1(1'b0), .CI(n2877), .O(n2874), .CO(n2875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i4 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i3  (.I0(\u_sensor_frame_count/cmos_fps_cnt[2] ), 
            .I1(1'b0), .CI(n602), .O(n2876), .CO(n2877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i3 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i28  (.I0(\u_sensor_frame_count/delay_cnt[27] ), 
            .I1(1'b0), .CI(n2880), .O(n2878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i28 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i27  (.I0(\u_sensor_frame_count/delay_cnt[26] ), 
            .I1(1'b0), .CI(n2882), .O(n2879), .CO(n2880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i27 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i26  (.I0(\u_sensor_frame_count/delay_cnt[25] ), 
            .I1(1'b0), .CI(n2884), .O(n2881), .CO(n2882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i26 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i25  (.I0(\u_sensor_frame_count/delay_cnt[24] ), 
            .I1(1'b0), .CI(n2886), .O(n2883), .CO(n2884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i25 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i24  (.I0(\u_sensor_frame_count/delay_cnt[23] ), 
            .I1(1'b0), .CI(n2888), .O(n2885), .CO(n2886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i24 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i23  (.I0(\u_sensor_frame_count/delay_cnt[22] ), 
            .I1(1'b0), .CI(n2890), .O(n2887), .CO(n2888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i23 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i22  (.I0(\u_sensor_frame_count/delay_cnt[21] ), 
            .I1(1'b0), .CI(n2892), .O(n2889), .CO(n2890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i22 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i21  (.I0(\u_sensor_frame_count/delay_cnt[20] ), 
            .I1(1'b0), .CI(n2909), .O(n2891), .CO(n2892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i21 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i20  (.I0(\u_sensor_frame_count/delay_cnt[19] ), 
            .I1(1'b0), .CI(n2911), .O(n2908), .CO(n2909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i20 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i19  (.I0(\u_sensor_frame_count/delay_cnt[18] ), 
            .I1(1'b0), .CI(n3042), .O(n2910), .CO(n2911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i19 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i2  (.I0(\u_lcd_driver/vcnt[1] ), .I1(\u_lcd_driver/vcnt[0] ), 
            .CI(1'b0), .O(n3039), .CO(n3040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i2 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i18  (.I0(\u_sensor_frame_count/delay_cnt[17] ), 
            .I1(1'b0), .CI(n3046), .O(n3041), .CO(n3042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i18 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i17  (.I0(\u_sensor_frame_count/delay_cnt[16] ), 
            .I1(1'b0), .CI(n3050), .O(n3045), .CO(n3046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i17 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_75/i2  (.I0(n371), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q_pinv ), 
            .CI(1'b0), .O(n3047), .CO(n3048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_0/add_75/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_75/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_sensor_frame_count/add_14/i16  (.I0(\u_sensor_frame_count/delay_cnt[15] ), 
            .I1(1'b0), .CI(n3054), .O(n3049), .CO(n3050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i16 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i15  (.I0(\u_sensor_frame_count/delay_cnt[14] ), 
            .I1(1'b0), .CI(n3056), .O(n3053), .CO(n3054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i15 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i14  (.I0(\u_sensor_frame_count/delay_cnt[13] ), 
            .I1(1'b0), .CI(n3061), .O(n3055), .CO(n3056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i14 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i13  (.I0(\u_sensor_frame_count/delay_cnt[12] ), 
            .I1(1'b0), .CI(n3063), .O(n3060), .CO(n3061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i13 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i12  (.I0(\u_sensor_frame_count/delay_cnt[11] ), 
            .I1(1'b0), .CI(n3076), .O(n3062), .CO(n3063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i12 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i11  (.I0(\u_sensor_frame_count/delay_cnt[10] ), 
            .I1(1'b0), .CI(n3078), .O(n3075), .CO(n3076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i11 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i10  (.I0(\u_sensor_frame_count/delay_cnt[9] ), 
            .I1(1'b0), .CI(n3080), .O(n3077), .CO(n3078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i10 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i9  (.I0(\u_sensor_frame_count/delay_cnt[8] ), 
            .I1(1'b0), .CI(n3082), .O(n3079), .CO(n3080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i9 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i8  (.I0(\u_sensor_frame_count/delay_cnt[7] ), 
            .I1(1'b0), .CI(n3084), .O(n3081), .CO(n3082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i8 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i7  (.I0(\u_sensor_frame_count/delay_cnt[6] ), 
            .I1(1'b0), .CI(n3086), .O(n3083), .CO(n3084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i7 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i6  (.I0(\u_sensor_frame_count/delay_cnt[5] ), 
            .I1(1'b0), .CI(n3088), .O(n3085), .CO(n3086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i6 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i5  (.I0(\u_sensor_frame_count/delay_cnt[4] ), 
            .I1(1'b0), .CI(n3090), .O(n3087), .CO(n3088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i5 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i4  (.I0(\u_sensor_frame_count/delay_cnt[3] ), 
            .I1(1'b0), .CI(n3092), .O(n3089), .CO(n3090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i4 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i3  (.I0(\u_sensor_frame_count/delay_cnt[2] ), 
            .I1(1'b0), .CI(n576), .O(n3091), .CO(n3092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i3 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i1  (.I0(\u_rgb2dvi/enc_0/acc[0] ), .I1(n3343), 
            .CI(1'b0), .O(n3203), .CO(n3204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i2  (.I0(n378), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q_pinv ), 
            .CI(n10604), .O(n3217), .CO(n3218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i12  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[11] ), 
            .I1(1'b0), .CI(n3221), .O(n3219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i12 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i11  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[10] ), 
            .I1(1'b0), .CI(n3223), .O(n3220), .CO(n3221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i11 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i10  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[9] ), 
            .I1(1'b0), .CI(n3225), .O(n3222), .CO(n3223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i10 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i9  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[8] ), 
            .I1(1'b0), .CI(n3227), .O(n3224), .CO(n3225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i9 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i8  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[7] ), 
            .I1(1'b0), .CI(n3229), .O(n3226), .CO(n3227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i8 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i7  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[6] ), 
            .I1(1'b0), .CI(n3231), .O(n3228), .CO(n3229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i7 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i6  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[5] ), 
            .I1(1'b0), .CI(n3233), .O(n3230), .CO(n3231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i6 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i5  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[4] ), 
            .I1(1'b0), .CI(n3235), .O(n3232), .CO(n3233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i5 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i4  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[3] ), 
            .I1(1'b0), .CI(n3237), .O(n3234), .CO(n3235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i4 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i3  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[2] ), 
            .I1(1'b0), .CI(n446), .O(n3236), .CO(n3237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i3 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i1  (.I0(\u_rgb2dvi/enc_1/acc[0] ), .I1(n3343), 
            .CI(1'b0), .O(n3282), .CO(n3283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i8  (.I0(\i2c_config_index[7] ), 
            .I1(1'b0), .CI(n3296), .O(n3294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i8 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i7  (.I0(\i2c_config_index[6] ), 
            .I1(1'b0), .CI(n3298), .O(n3295), .CO(n3296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i7 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i6  (.I0(\i2c_config_index[5] ), 
            .I1(1'b0), .CI(n3300), .O(n3297), .CO(n3298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i6 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i5  (.I0(\i2c_config_index[4] ), 
            .I1(1'b0), .CI(n3302), .O(n3299), .CO(n3300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i5 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i4  (.I0(\i2c_config_index[3] ), 
            .I1(1'b0), .CI(n3304), .O(n3301), .CO(n3302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i4 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i3  (.I0(\i2c_config_index[2] ), 
            .I1(1'b0), .CI(n232), .O(n3303), .CO(n3304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i3 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i16  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15] ), 
            .I1(1'b0), .CI(n3307), .O(n3305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i16 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i15  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14] ), 
            .I1(1'b0), .CI(n3318), .O(n3306), .CO(n3307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i15 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i14  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13] ), 
            .I1(1'b0), .CI(n3320), .O(n3317), .CO(n3318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i14 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i13  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), 
            .I1(1'b0), .CI(n3322), .O(n3319), .CO(n3320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i13 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i12  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] ), 
            .I1(1'b0), .CI(n3324), .O(n3321), .CO(n3322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i12 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i11  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), 
            .I1(1'b0), .CI(n3330), .O(n3323), .CO(n3324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i11 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i10  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), 
            .I1(1'b0), .CI(n3332), .O(n3329), .CO(n3330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i10 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i9  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] ), 
            .I1(1'b0), .CI(n3334), .O(n3331), .CO(n3332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i9 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i8  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), 
            .I1(1'b0), .CI(n3336), .O(n3333), .CO(n3334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i8 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i7  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] ), 
            .I1(1'b0), .CI(n3338), .O(n3335), .CO(n3336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i7 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i6  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] ), 
            .I1(1'b0), .CI(n3342), .O(n3337), .CO(n3338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i6 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i1  (.I0(\u_rgb2dvi/enc_2/acc[0] ), .I1(n3343), 
            .CI(1'b0), .O(n3339), .CO(n3340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i5  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4] ), 
            .I1(1'b0), .CI(n3347), .O(n3341), .CO(n3342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i5 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/sub_50/add_2/i1  (.I0(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q ), .CI(n10605), .O(n3343), 
            .CO(n10606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_2/sub_50/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/sub_50/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i4  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3] ), 
            .I1(1'b0), .CI(n3349), .O(n3346), .CO(n3347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i4 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i3  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2] ), 
            .I1(1'b0), .CI(n229), .O(n3348), .CO(n3349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i3 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i20  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19] ), 
            .I1(1'b0), .CI(n3353), .O(n3351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i20 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i19  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18] ), 
            .I1(1'b0), .CI(n3355), .O(n3352), .CO(n3353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i19 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i18  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17] ), 
            .I1(1'b0), .CI(n3357), .O(n3354), .CO(n3355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i18 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i17  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16] ), 
            .I1(1'b0), .CI(n3359), .O(n3356), .CO(n3357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i17 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i16  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15] ), 
            .I1(1'b0), .CI(n3361), .O(n3358), .CO(n3359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i16 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i15  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14] ), 
            .I1(1'b0), .CI(n3363), .O(n3360), .CO(n3361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i15 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i14  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13] ), 
            .I1(1'b0), .CI(n3365), .O(n3362), .CO(n3363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i14 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i13  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12] ), 
            .I1(1'b0), .CI(n3367), .O(n3364), .CO(n3365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i13 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i12  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11] ), 
            .I1(1'b0), .CI(n3369), .O(n3366), .CO(n3367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i12 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i11  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10] ), 
            .I1(1'b0), .CI(n3379), .O(n3368), .CO(n3369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i11 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i10  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9] ), 
            .I1(1'b0), .CI(n3381), .O(n3378), .CO(n3379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i10 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i9  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8] ), 
            .I1(1'b0), .CI(n3383), .O(n3380), .CO(n3381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i9 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i8  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7] ), 
            .I1(1'b0), .CI(n3385), .O(n3382), .CO(n3383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i8 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i7  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6] ), 
            .I1(1'b0), .CI(n3387), .O(n3384), .CO(n3385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i7 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i6  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5] ), 
            .I1(1'b0), .CI(n3389), .O(n3386), .CO(n3387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i6 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i5  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4] ), 
            .I1(1'b0), .CI(n3391), .O(n3388), .CO(n3389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i5 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i4  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3] ), 
            .I1(1'b0), .CI(n3393), .O(n3390), .CO(n3391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i4 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i3  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2] ), 
            .I1(1'b0), .CI(n206), .O(n3392), .CO(n3393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i3 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] ), 
            .I1(1'b1), .CI(n3400), .O(n3398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] ), 
            .I1(1'b1), .CI(n3402), .O(n3399), .CO(n3400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] ), 
            .I1(1'b1), .CI(n3404), .O(n3401), .CO(n3402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] ), 
            .I1(1'b1), .CI(n3406), .O(n3403), .CO(n3404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] ), 
            .I1(1'b1), .CI(n3408), .O(n3405), .CO(n3406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] ), 
            .I1(1'b1), .CI(n3410), .O(n3407), .CO(n3408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] ), 
            .I1(1'b1), .CI(n3412), .O(n3409), .CO(n3410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] ), 
            .I1(1'b1), .CI(n3414), .O(n3411), .CO(n3412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] ), 
            .I1(1'b1), .CI(n3416), .O(n3413), .CO(n3414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] ), 
            .I1(1'b1), .CI(n3418), .O(n3415), .CO(n3416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] ), 
            .I1(1'b1), .CI(n3420), .O(n3417), .CO(n3418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] ), 
            .I1(1'b1), .CI(n3422), .O(n3419), .CO(n3420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] ), 
            .I1(1'b1), .CI(n3424), .O(n3421), .CO(n3422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] ), 
            .I1(1'b1), .CI(n3426), .O(n3423), .CO(n3424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] ), 
            .I1(1'b1), .CI(n3428), .O(n3425), .CO(n3426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] ), 
            .I1(1'b1), .CI(n3430), .O(n3427), .CO(n3428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] ), 
            .I1(1'b1), .CI(n3432), .O(n3429), .CO(n3430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] ), 
            .I1(1'b1), .CI(n3434), .O(n3431), .CO(n3432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] ), 
            .I1(1'b1), .CI(n187), .O(n3433), .CO(n3434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i8  (.I0(\PowerOnResetCnt[7] ), .I1(1'b0), .CI(n3438), 
            .O(n3436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i8 .I0_POLARITY = 1'b1;
    defparam \add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i7  (.I0(\PowerOnResetCnt[6] ), .I1(1'b0), .CI(n3440), 
            .O(n3437), .CO(n3438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i7 .I0_POLARITY = 1'b1;
    defparam \add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i6  (.I0(\PowerOnResetCnt[5] ), .I1(1'b0), .CI(n3442), 
            .O(n3439), .CO(n3440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i6 .I0_POLARITY = 1'b1;
    defparam \add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i5  (.I0(\PowerOnResetCnt[4] ), .I1(1'b0), .CI(n4985), 
            .O(n3441), .CO(n3442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i5 .I0_POLARITY = 1'b1;
    defparam \add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i4  (.I0(\PowerOnResetCnt[3] ), .I1(1'b0), .CI(n4987), 
            .O(n4984), .CO(n4985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i4 .I0_POLARITY = 1'b1;
    defparam \add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i3  (.I0(\PowerOnResetCnt[2] ), .I1(1'b0), .CI(n4989), 
            .O(n4986), .CO(n4987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i3 .I0_POLARITY = 1'b1;
    defparam \add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i2  (.I0(\PowerOnResetCnt[1] ), .I1(1'b0), .CI(n4991), 
            .O(n4988), .CO(n4989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i2 .I0_POLARITY = 1'b1;
    defparam \add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i1  (.I0(\PowerOnResetCnt[0] ), .I1(\reduce_nand_9/n7 ), 
            .CI(1'b0), .O(n4990), .CO(n4991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i1 .I0_POLARITY = 1'b1;
    defparam \add_10/i1 .I1_POLARITY = 1'b0;
    EFX_LUT4 \edb_top_inst/LUT__2678  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/edb_user_dr[62] ), .I2(\edb_top_inst/la0/crc_data_out[13] ), 
            .I3(\edb_top_inst/edb_user_dr[63] ), .O(\edb_top_inst/n1731 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2678 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2679  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/edb_user_dr[57] ), .I2(\edb_top_inst/la0/crc_data_out[14] ), 
            .I3(\edb_top_inst/edb_user_dr[64] ), .O(\edb_top_inst/n1732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2679 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2680  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/edb_user_dr[58] ), .I2(\edb_top_inst/la0/crc_data_out[9] ), 
            .I3(\edb_top_inst/edb_user_dr[59] ), .O(\edb_top_inst/n1733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2680 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2681  (.I0(\edb_top_inst/n1730 ), .I1(\edb_top_inst/n1731 ), 
            .I2(\edb_top_inst/n1732 ), .I3(\edb_top_inst/n1733 ), .O(\edb_top_inst/n1734 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2681 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__2682  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/edb_user_dr[52] ), .I2(\edb_top_inst/la0/crc_data_out[3] ), 
            .I3(\edb_top_inst/edb_user_dr[53] ), .O(\edb_top_inst/n1735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2682 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2683  (.I0(\edb_top_inst/la0/crc_data_out[0] ), 
            .I1(\edb_top_inst/edb_user_dr[50] ), .I2(\edb_top_inst/la0/crc_data_out[1] ), 
            .I3(\edb_top_inst/edb_user_dr[51] ), .O(\edb_top_inst/n1736 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2683 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2684  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/edb_user_dr[54] ), .I2(\edb_top_inst/la0/crc_data_out[5] ), 
            .I3(\edb_top_inst/edb_user_dr[55] ), .O(\edb_top_inst/n1737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2684 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2685  (.I0(\edb_top_inst/la0/crc_data_out[6] ), 
            .I1(\edb_top_inst/edb_user_dr[56] ), .I2(\edb_top_inst/la0/crc_data_out[15] ), 
            .I3(\edb_top_inst/edb_user_dr[65] ), .O(\edb_top_inst/n1738 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2685 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2686  (.I0(\edb_top_inst/n1735 ), .I1(\edb_top_inst/n1736 ), 
            .I2(\edb_top_inst/n1737 ), .I3(\edb_top_inst/n1738 ), .O(\edb_top_inst/n1739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2686 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__2687  (.I0(\edb_top_inst/la0/crc_data_out[16] ), 
            .I1(\edb_top_inst/edb_user_dr[66] ), .I2(\edb_top_inst/la0/crc_data_out[23] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n1740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2687 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2688  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/edb_user_dr[67] ), .I2(\edb_top_inst/la0/crc_data_out[18] ), 
            .I3(\edb_top_inst/edb_user_dr[68] ), .O(\edb_top_inst/n1741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2688 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2689  (.I0(\edb_top_inst/la0/crc_data_out[21] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/la0/crc_data_out[22] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/n1742 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2689 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2690  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/edb_user_dr[69] ), .I2(\edb_top_inst/la0/crc_data_out[20] ), 
            .I3(\edb_top_inst/edb_user_dr[70] ), .O(\edb_top_inst/n1743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2690 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2691  (.I0(\edb_top_inst/n1740 ), .I1(\edb_top_inst/n1741 ), 
            .I2(\edb_top_inst/n1742 ), .I3(\edb_top_inst/n1743 ), .O(\edb_top_inst/n1744 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2691 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__2692  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/edb_user_dr[79] ), .I2(\edb_top_inst/la0/crc_data_out[30] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n1745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2692 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2693  (.I0(\edb_top_inst/la0/crc_data_out[25] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/la0/crc_data_out[26] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n1746 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2693 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2694  (.I0(\edb_top_inst/la0/crc_data_out[27] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/la0/crc_data_out[28] ), 
            .I3(\edb_top_inst/edb_user_dr[78] ), .O(\edb_top_inst/n1747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2694 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2695  (.I0(\edb_top_inst/la0/crc_data_out[24] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/la0/crc_data_out[31] ), 
            .I3(\edb_top_inst/edb_user_dr[81] ), .O(\edb_top_inst/n1748 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2695 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__2696  (.I0(\edb_top_inst/n1745 ), .I1(\edb_top_inst/n1746 ), 
            .I2(\edb_top_inst/n1747 ), .I3(\edb_top_inst/n1748 ), .O(\edb_top_inst/n1749 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2696 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__2697  (.I0(\edb_top_inst/n1734 ), .I1(\edb_top_inst/n1739 ), 
            .I2(\edb_top_inst/n1744 ), .I3(\edb_top_inst/n1749 ), .O(\edb_top_inst/n1750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2697 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__2698  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/la0/bit_count[2] ), 
            .O(\edb_top_inst/n1751 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2698 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__2699  (.I0(\edb_top_inst/la0/bit_count[3] ), 
            .I1(\edb_top_inst/la0/bit_count[4] ), .I2(\edb_top_inst/la0/bit_count[5] ), 
            .O(\edb_top_inst/n1752 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2699 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__2700  (.I0(\edb_top_inst/n1752 ), .I1(\edb_top_inst/n1751 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n1753 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2700 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__2701  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/n1753 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n1754 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2701 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__2702  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/n1754 ), .O(\edb_top_inst/n1755 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2702 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2703  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n1756 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2703 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2704  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/n1755 ), .I2(\edb_top_inst/n1756 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n1757 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2704 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__2705  (.I0(\edb_top_inst/n1750 ), .I1(\edb_top_inst/la0/biu_ready ), 
            .I2(\edb_top_inst/n1757 ), .O(\edb_top_inst/n1758 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2705 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2706  (.I0(\edb_top_inst/la0/crc_data_out[0] ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), .I2(\edb_top_inst/n1757 ), 
            .O(\edb_top_inst/n1759 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2706 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2707  (.I0(\edb_top_inst/n1754 ), .I1(\edb_top_inst/la0/module_state[1] ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n1760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2707 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__2708  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n1761 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2708 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2709  (.I0(\edb_top_inst/n1760 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/n1761 ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n1762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2709 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__2710  (.I0(\edb_top_inst/debug_hub_inst/module_id_reg[1] ), 
            .I1(\edb_top_inst/debug_hub_inst/module_id_reg[2] ), .I2(\edb_top_inst/debug_hub_inst/module_id_reg[3] ), 
            .I3(\edb_top_inst/debug_hub_inst/module_id_reg[0] ), .O(\edb_top_inst/n1763 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2710 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__2711  (.I0(\edb_top_inst/n1759 ), .I1(\edb_top_inst/n1758 ), 
            .I2(\edb_top_inst/n1762 ), .I3(\edb_top_inst/n1763 ), .O(jtag_inst1_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2711 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__2712  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[40] ), .O(\edb_top_inst/la0/n1317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2712 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2713  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/edb_user_dr[67] ), .I2(\edb_top_inst/edb_user_dr[68] ), 
            .I3(\edb_top_inst/edb_user_dr[69] ), .O(\edb_top_inst/n1764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2713 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2714  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .O(\edb_top_inst/n1765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2714 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2715  (.I0(\edb_top_inst/n1764 ), .I1(\edb_top_inst/n1765 ), 
            .O(\edb_top_inst/n1766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2715 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__2716  (.I0(\edb_top_inst/edb_user_dr[74] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/edb_user_dr[76] ), 
            .I3(\edb_top_inst/edb_user_dr[79] ), .O(\edb_top_inst/n1767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2716 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2717  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .I2(\edb_top_inst/n1756 ), 
            .O(\edb_top_inst/n1768 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2717 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__2718  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(jtag_inst1_UPDATE), .O(\edb_top_inst/n1769 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2718 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2719  (.I0(\edb_top_inst/n1763 ), .I1(\edb_top_inst/n1768 ), 
            .I2(\edb_top_inst/n1769 ), .O(\edb_top_inst/n1770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2719 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__2720  (.I0(\edb_top_inst/edb_user_dr[78] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/edb_user_dr[80] ), 
            .I3(\edb_top_inst/n1770 ), .O(\edb_top_inst/la0/regsel_ld_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2720 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__2721  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[73] ), .I2(\edb_top_inst/n1767 ), 
            .I3(\edb_top_inst/la0/regsel_ld_en ), .O(\edb_top_inst/n1771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2721 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__2722  (.I0(\edb_top_inst/edb_user_dr[71] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/n1771 ), 
            .O(\edb_top_inst/n1772 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2722 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__2723  (.I0(\edb_top_inst/n1772 ), .I1(\edb_top_inst/n1766 ), 
            .I2(\edb_top_inst/la0/la_soft_reset_in ), .O(\edb_top_inst/ceg_net5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2723 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__2724  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/n1766 ), .I2(\edb_top_inst/n1772 ), .O(\edb_top_inst/la0/n6737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2724 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__2725  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[41] ), .O(\edb_top_inst/la0/n1318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2725 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2726  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[42] ), .O(\edb_top_inst/la0/n1319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2726 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2727  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/edb_user_dr[64] ), .I2(\edb_top_inst/n1764 ), 
            .I3(\edb_top_inst/n1772 ), .O(\edb_top_inst/la0/n1373 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2727 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__2728  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n1764 ), 
            .I3(\edb_top_inst/n1772 ), .O(\edb_top_inst/la0/n1890 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2728 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__2729  (.I0(\edb_top_inst/edb_user_dr[67] ), 
            .I1(\edb_top_inst/edb_user_dr[68] ), .I2(\edb_top_inst/edb_user_dr[63] ), 
            .I3(\edb_top_inst/edb_user_dr[66] ), .O(\edb_top_inst/n1773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2729 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__2730  (.I0(\edb_top_inst/edb_user_dr[69] ), 
            .I1(\edb_top_inst/n1765 ), .I2(\edb_top_inst/n1772 ), .I3(\edb_top_inst/n1773 ), 
            .O(\edb_top_inst/la0/n1942 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2730 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__2731  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(\edb_top_inst/la0/address_counter[9] ), .I2(\edb_top_inst/la0/address_counter[10] ), 
            .I3(\edb_top_inst/la0/address_counter[11] ), .O(\edb_top_inst/n1774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2731 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2732  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/la0/address_counter[12] ), .I2(\edb_top_inst/la0/address_counter[13] ), 
            .I3(\edb_top_inst/la0/address_counter[14] ), .O(\edb_top_inst/n1775 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2732 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2733  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(\edb_top_inst/la0/address_counter[5] ), .I2(\edb_top_inst/la0/address_counter[6] ), 
            .I3(\edb_top_inst/la0/address_counter[7] ), .O(\edb_top_inst/n1776 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2733 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2734  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/la0/address_counter[1] ), .I2(\edb_top_inst/la0/address_counter[2] ), 
            .O(\edb_top_inst/n1777 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2734 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__2735  (.I0(\edb_top_inst/n1774 ), .I1(\edb_top_inst/n1775 ), 
            .I2(\edb_top_inst/n1776 ), .I3(\edb_top_inst/n1777 ), .O(\edb_top_inst/n1778 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2735 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__2736  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n34 ), 
            .I2(\edb_top_inst/edb_user_dr[45] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2736 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2737  (.I0(\edb_top_inst/edb_user_dr[77] ), 
            .I1(\edb_top_inst/edb_user_dr[78] ), .I2(\edb_top_inst/edb_user_dr[79] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n1779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2737 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__2738  (.I0(\edb_top_inst/n1779 ), .I1(\edb_top_inst/n1768 ), 
            .I2(\edb_top_inst/n1769 ), .I3(\edb_top_inst/n1763 ), .O(\edb_top_inst/n1780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2738 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__2739  (.I0(\edb_top_inst/la0/word_count[6] ), 
            .I1(\edb_top_inst/la0/word_count[7] ), .I2(\edb_top_inst/la0/word_count[8] ), 
            .I3(\edb_top_inst/la0/word_count[9] ), .O(\edb_top_inst/n1781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2739 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2740  (.I0(\edb_top_inst/la0/word_count[1] ), 
            .I1(\edb_top_inst/la0/word_count[2] ), .I2(\edb_top_inst/la0/word_count[3] ), 
            .O(\edb_top_inst/n1782 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2740 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__2741  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/la0/word_count[13] ), .I2(\edb_top_inst/la0/word_count[14] ), 
            .I3(\edb_top_inst/la0/word_count[15] ), .O(\edb_top_inst/n1783 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2741 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2742  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/la0/word_count[10] ), 
            .I3(\edb_top_inst/la0/word_count[11] ), .O(\edb_top_inst/n1784 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2742 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2743  (.I0(\edb_top_inst/n1781 ), .I1(\edb_top_inst/n1782 ), 
            .I2(\edb_top_inst/n1783 ), .I3(\edb_top_inst/n1784 ), .O(\edb_top_inst/n1785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2743 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__2744  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/n1785 ), .O(\edb_top_inst/n1786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2744 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2745  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n1787 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2745 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2746  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n1788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2746 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__2747  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n1789 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2747 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__2748  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/la0/bit_count[2] ), 
            .I3(\edb_top_inst/n1789 ), .O(\edb_top_inst/n1790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe7f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2748 .LUTMASK = 16'hfe7f;
    EFX_LUT4 \edb_top_inst/LUT__2749  (.I0(\edb_top_inst/la0/opcode[3] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/n1708 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2749 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__2750  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n1705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2750 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__2751  (.I0(\edb_top_inst/n1708 ), .I1(\edb_top_inst/la0/bit_count[5] ), 
            .I2(\edb_top_inst/n1705 ), .I3(\edb_top_inst/la0/bit_count[4] ), 
            .O(\edb_top_inst/n1791 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2751 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__2752  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n1792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2752 .LUTMASK = 16'hfe3f;
    EFX_LUT4 \edb_top_inst/LUT__2753  (.I0(\edb_top_inst/n1790 ), .I1(\edb_top_inst/n1791 ), 
            .I2(\edb_top_inst/la0/bit_count[3] ), .I3(\edb_top_inst/n1792 ), 
            .O(\edb_top_inst/n1793 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2753 .LUTMASK = 16'h0110;
    EFX_LUT4 \edb_top_inst/LUT__2754  (.I0(\edb_top_inst/n1786 ), .I1(\edb_top_inst/n1787 ), 
            .I2(\edb_top_inst/n1788 ), .I3(\edb_top_inst/n1793 ), .O(\edb_top_inst/n1794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5333, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2754 .LUTMASK = 16'h5333;
    EFX_LUT4 \edb_top_inst/LUT__2755  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/la0/biu_ready ), .O(\edb_top_inst/n1795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2755 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__2756  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .I3(\edb_top_inst/la0/word_count[3] ), .O(\edb_top_inst/n1796 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2756 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2757  (.I0(\edb_top_inst/n1781 ), .I1(\edb_top_inst/n1783 ), 
            .I2(\edb_top_inst/n1784 ), .I3(\edb_top_inst/n1796 ), .O(\edb_top_inst/n1797 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2757 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__2758  (.I0(\edb_top_inst/n1797 ), .I1(\edb_top_inst/n1761 ), 
            .O(\edb_top_inst/n1798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2758 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2759  (.I0(\edb_top_inst/n1795 ), .I1(\edb_top_inst/n1785 ), 
            .I2(\edb_top_inst/n1798 ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n1799 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2759 .LUTMASK = 16'h000d;
    EFX_LUT4 \edb_top_inst/LUT__2760  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/n1756 ), .O(\edb_top_inst/n1800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2760 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2761  (.I0(\edb_top_inst/n1799 ), .I1(\edb_top_inst/n1794 ), 
            .I2(\edb_top_inst/n1800 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n1801 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2761 .LUTMASK = 16'h0fbb;
    EFX_LUT4 \edb_top_inst/LUT__2762  (.I0(\edb_top_inst/n1780 ), .I1(\edb_top_inst/n1801 ), 
            .O(\edb_top_inst/la0/addr_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2762 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__2763  (.I0(\edb_top_inst/la0/opcode[1] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/n969 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2763 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__2764  (.I0(\edb_top_inst/n1779 ), .I1(\edb_top_inst/n1770 ), 
            .O(\edb_top_inst/la0/op_reg_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2764 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2765  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/n1795 ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n1802 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2765 .LUTMASK = 16'h00f8;
    EFX_LUT4 \edb_top_inst/LUT__2766  (.I0(\edb_top_inst/n1780 ), .I1(\edb_top_inst/la0/module_state[3] ), 
            .I2(\edb_top_inst/n1800 ), .O(\edb_top_inst/n1803 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2766 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__2767  (.I0(\edb_top_inst/n1788 ), .I1(\edb_top_inst/n1793 ), 
            .I2(\edb_top_inst/n1787 ), .O(\edb_top_inst/n1804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2767 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__2768  (.I0(\edb_top_inst/n1803 ), .I1(\edb_top_inst/n1802 ), 
            .I2(\edb_top_inst/n1804 ), .O(\edb_top_inst/n1805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2768 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__2769  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/n1805 ), .O(\edb_top_inst/la0/n2166 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2769 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2770  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .I2(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n1806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2770 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__2771  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n1807 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2771 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2772  (.I0(\edb_top_inst/n1807 ), .I1(\edb_top_inst/edb_user_dr[81] ), 
            .I2(\edb_top_inst/n1763 ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n1808 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2772 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__2773  (.I0(\edb_top_inst/n1808 ), .I1(\edb_top_inst/n1755 ), 
            .I2(\edb_top_inst/n1787 ), .O(\edb_top_inst/n1809 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2773 .LUTMASK = 16'h6060;
    EFX_LUT4 \edb_top_inst/LUT__2774  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n1809 ), .O(\edb_top_inst/n1810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2774 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2775  (.I0(\edb_top_inst/n1802 ), .I1(\edb_top_inst/n1794 ), 
            .I2(\edb_top_inst/n1806 ), .I3(\edb_top_inst/n1810 ), .O(\edb_top_inst/ceg_net26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2775 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__2776  (.I0(\edb_top_inst/edb_user_dr[29] ), 
            .I1(\edb_top_inst/la0/word_count[0] ), .I2(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_word_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2776 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__2777  (.I0(\edb_top_inst/n1793 ), .I1(\edb_top_inst/n1797 ), 
            .O(\edb_top_inst/n1811 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2777 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__2778  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n1812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2778 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2779  (.I0(\edb_top_inst/n1811 ), .I1(\edb_top_inst/n1812 ), 
            .I2(\edb_top_inst/n1808 ), .I3(\edb_top_inst/n1787 ), .O(\edb_top_inst/n1813 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2779 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__2780  (.I0(jtag_inst1_CAPTURE), .I1(\edb_top_inst/n1763 ), 
            .O(\edb_top_inst/n1814 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2780 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__2781  (.I0(\edb_top_inst/n1797 ), .I1(\edb_top_inst/n1814 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n1815 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2781 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__2782  (.I0(\edb_top_inst/n1811 ), .I1(\edb_top_inst/n1807 ), 
            .I2(\edb_top_inst/n1815 ), .O(\edb_top_inst/n1816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2782 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__2783  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .I2(jtag_inst1_UPDATE), 
            .O(\edb_top_inst/n1817 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2783 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__2784  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .I2(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n1818 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2784 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__2785  (.I0(\edb_top_inst/n1814 ), .I1(\edb_top_inst/n1817 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/n1818 ), 
            .O(\edb_top_inst/n1819 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2785 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__2786  (.I0(\edb_top_inst/n1756 ), .I1(\edb_top_inst/n1797 ), 
            .I2(\edb_top_inst/n1754 ), .I3(\edb_top_inst/n1819 ), .O(\edb_top_inst/n1820 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2786 .LUTMASK = 16'h008f;
    EFX_LUT4 \edb_top_inst/LUT__2787  (.I0(\edb_top_inst/n1816 ), .I1(\edb_top_inst/n1813 ), 
            .I2(\edb_top_inst/n1780 ), .I3(\edb_top_inst/n1820 ), .O(\edb_top_inst/la0/module_next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2787 .LUTMASK = 16'hf4ff;
    EFX_LUT4 \edb_top_inst/LUT__2788  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .I2(\edb_top_inst/la0/module_next_state[0] ), 
            .I3(\edb_top_inst/n1805 ), .O(\edb_top_inst/la0/word_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2788 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__2789  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n1821 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hec07, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2789 .LUTMASK = 16'hec07;
    EFX_LUT4 \edb_top_inst/LUT__2790  (.I0(\edb_top_inst/n1821 ), .I1(\edb_top_inst/la0/la_trig_mask[0] ), 
            .I2(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1822 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2790 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__2791  (.I0(\edb_top_inst/la0/internal_register_select[10] ), 
            .I1(\edb_top_inst/la0/internal_register_select[11] ), .O(\edb_top_inst/n1823 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2791 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2792  (.I0(\edb_top_inst/la0/internal_register_select[1] ), 
            .I1(\edb_top_inst/la0/internal_register_select[2] ), .I2(\edb_top_inst/la0/internal_register_select[4] ), 
            .I3(\edb_top_inst/la0/internal_register_select[5] ), .O(\edb_top_inst/n1824 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2792 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2793  (.I0(\edb_top_inst/la0/internal_register_select[6] ), 
            .I1(\edb_top_inst/la0/internal_register_select[7] ), .I2(\edb_top_inst/la0/internal_register_select[8] ), 
            .I3(\edb_top_inst/la0/internal_register_select[9] ), .O(\edb_top_inst/n1825 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2793 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__2794  (.I0(\edb_top_inst/la0/internal_register_select[12] ), 
            .I1(\edb_top_inst/n1823 ), .I2(\edb_top_inst/n1824 ), .I3(\edb_top_inst/n1825 ), 
            .O(\edb_top_inst/n1826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2794 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__2795  (.I0(\edb_top_inst/n1802 ), .I1(\edb_top_inst/n1826 ), 
            .O(\edb_top_inst/n1827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2795 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2796  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/n1827 ), .O(\edb_top_inst/n1828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2796 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2797  (.I0(\edb_top_inst/n1822 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_from_biu[0] ), .I3(\edb_top_inst/n1802 ), 
            .O(\edb_top_inst/n1829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2797 .LUTMASK = 16'h0bbb;
    EFX_LUT4 \edb_top_inst/LUT__2798  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n1756 ), .I2(\edb_top_inst/n1814 ), .I3(\edb_top_inst/n1802 ), 
            .O(\edb_top_inst/n1830 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2798 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__2799  (.I0(\edb_top_inst/n1756 ), .I1(\edb_top_inst/n1793 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/n1830 ), 
            .O(\edb_top_inst/n1831 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2799 .LUTMASK = 16'h008f;
    EFX_LUT4 \edb_top_inst/LUT__2800  (.I0(\edb_top_inst/n1829 ), .I1(\edb_top_inst/la0/data_out_shift_reg[1] ), 
            .I2(\edb_top_inst/n1831 ), .O(\edb_top_inst/la0/n2443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2800 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__2801  (.I0(\edb_top_inst/n1763 ), .I1(jtag_inst1_SHIFT), 
            .I2(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n1832 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2801 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__2802  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n1832 ), .I2(\edb_top_inst/n1756 ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/ceg_net14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2802 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__2803  (.I0(jtag_inst1_RESET), .I1(\edb_top_inst/la0/la_soft_reset_in ), 
            .O(\edb_top_inst/la0/n2730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2803 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__2804  (.I0(\edb_top_inst/edb_user_dr[72] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/n1766 ), 
            .I3(\edb_top_inst/n1771 ), .O(\edb_top_inst/la0/n2743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2804 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__2805  (.I0(\edb_top_inst/edb_user_dr[71] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/n1766 ), 
            .I3(\edb_top_inst/n1771 ), .O(\edb_top_inst/la0/n3576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2805 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__2806  (.I0(\edb_top_inst/edb_user_dr[71] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/n1771 ), 
            .O(\edb_top_inst/n1833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2806 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__2807  (.I0(\edb_top_inst/n1766 ), .I1(\edb_top_inst/n1833 ), 
            .O(\edb_top_inst/la0/n4465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2807 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__2808  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/edb_user_dr[64] ), .I2(\edb_top_inst/n1764 ), 
            .I3(\edb_top_inst/n1833 ), .O(\edb_top_inst/la0/n4480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2808 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__2809  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n1764 ), 
            .I3(\edb_top_inst/n1833 ), .O(\edb_top_inst/la0/n4678 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2809 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__2810  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n833 ), 
            .I2(\edb_top_inst/edb_user_dr[46] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2810 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2811  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n831 ), 
            .I2(\edb_top_inst/edb_user_dr[47] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2811 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2812  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n829 ), 
            .I2(\edb_top_inst/edb_user_dr[48] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2812 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2813  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n827 ), 
            .I2(\edb_top_inst/edb_user_dr[49] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2813 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2814  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n825 ), 
            .I2(\edb_top_inst/edb_user_dr[50] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2814 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2815  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n823 ), 
            .I2(\edb_top_inst/edb_user_dr[51] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2815 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2816  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n821 ), 
            .I2(\edb_top_inst/edb_user_dr[52] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2816 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2817  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n819 ), 
            .I2(\edb_top_inst/edb_user_dr[53] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2817 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2818  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n817 ), 
            .I2(\edb_top_inst/edb_user_dr[54] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2818 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2819  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n815 ), 
            .I2(\edb_top_inst/edb_user_dr[55] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2819 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2820  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n813 ), 
            .I2(\edb_top_inst/edb_user_dr[56] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2820 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2821  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n811 ), 
            .I2(\edb_top_inst/edb_user_dr[57] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2821 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2822  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n809 ), 
            .I2(\edb_top_inst/edb_user_dr[58] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2822 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2823  (.I0(\edb_top_inst/n1778 ), .I1(\edb_top_inst/n807 ), 
            .I2(\edb_top_inst/edb_user_dr[59] ), .I3(\edb_top_inst/n1768 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2823 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__2824  (.I0(\edb_top_inst/n805 ), .I1(\edb_top_inst/la0/address_counter[15] ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2824 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2825  (.I0(\edb_top_inst/n1834 ), .I1(\edb_top_inst/edb_user_dr[60] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2825 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2826  (.I0(\edb_top_inst/n867 ), .I1(\edb_top_inst/n803 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1835 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2826 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2827  (.I0(\edb_top_inst/n1835 ), .I1(\edb_top_inst/edb_user_dr[61] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2827 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2828  (.I0(\edb_top_inst/n865 ), .I1(\edb_top_inst/n801 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2828 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2829  (.I0(\edb_top_inst/n1836 ), .I1(\edb_top_inst/edb_user_dr[62] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2829 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2830  (.I0(\edb_top_inst/n863 ), .I1(\edb_top_inst/n799 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1837 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2830 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2831  (.I0(\edb_top_inst/n1837 ), .I1(\edb_top_inst/edb_user_dr[63] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2831 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2832  (.I0(\edb_top_inst/n861 ), .I1(\edb_top_inst/n797 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2832 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2833  (.I0(\edb_top_inst/n1838 ), .I1(\edb_top_inst/edb_user_dr[64] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2833 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2834  (.I0(\edb_top_inst/n856 ), .I1(\edb_top_inst/n795 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2834 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2835  (.I0(\edb_top_inst/n1839 ), .I1(\edb_top_inst/edb_user_dr[65] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2835 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2836  (.I0(\edb_top_inst/n854 ), .I1(\edb_top_inst/n793 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2836 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2837  (.I0(\edb_top_inst/n1840 ), .I1(\edb_top_inst/edb_user_dr[66] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2837 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2838  (.I0(\edb_top_inst/n852 ), .I1(\edb_top_inst/n791 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2838 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2839  (.I0(\edb_top_inst/n1841 ), .I1(\edb_top_inst/edb_user_dr[67] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2839 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2840  (.I0(\edb_top_inst/n850 ), .I1(\edb_top_inst/n789 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2840 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2841  (.I0(\edb_top_inst/n1842 ), .I1(\edb_top_inst/edb_user_dr[68] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2841 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2842  (.I0(\edb_top_inst/n848 ), .I1(\edb_top_inst/n787 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2842 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2843  (.I0(\edb_top_inst/n1843 ), .I1(\edb_top_inst/edb_user_dr[69] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2843 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2844  (.I0(\edb_top_inst/n846 ), .I1(\edb_top_inst/n785 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2844 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2845  (.I0(\edb_top_inst/n1844 ), .I1(\edb_top_inst/edb_user_dr[70] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2845 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2846  (.I0(\edb_top_inst/n844 ), .I1(\edb_top_inst/n783 ), 
            .I2(\edb_top_inst/n1778 ), .O(\edb_top_inst/n1845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2846 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2847  (.I0(\edb_top_inst/n1845 ), .I1(\edb_top_inst/edb_user_dr[71] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_addr_counter[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2847 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2858  (.I0(\edb_top_inst/n1805 ), .I1(\edb_top_inst/n36 ), 
            .O(\edb_top_inst/la0/n2165 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2858 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2859  (.I0(\edb_top_inst/n1805 ), .I1(\edb_top_inst/n772 ), 
            .O(\edb_top_inst/la0/n2164 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2859 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2860  (.I0(\edb_top_inst/n1805 ), .I1(\edb_top_inst/n770 ), 
            .O(\edb_top_inst/la0/n2163 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2860 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2861  (.I0(\edb_top_inst/n1805 ), .I1(\edb_top_inst/n768 ), 
            .O(\edb_top_inst/la0/n2162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2861 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2862  (.I0(\edb_top_inst/n1805 ), .I1(\edb_top_inst/n767 ), 
            .O(\edb_top_inst/la0/n2161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2862 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2863  (.I0(\edb_top_inst/edb_user_dr[30] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[0] ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2863 .LUTMASK = 16'haac3;
    EFX_LUT4 \edb_top_inst/LUT__2864  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .O(\edb_top_inst/n1851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2864 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2865  (.I0(\edb_top_inst/edb_user_dr[31] ), 
            .I1(\edb_top_inst/la0/word_count[2] ), .I2(\edb_top_inst/n1851 ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2865 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__2866  (.I0(\edb_top_inst/la0/word_count[2] ), 
            .I1(\edb_top_inst/n1851 ), .I2(\edb_top_inst/la0/word_count[3] ), 
            .O(\edb_top_inst/n1852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2866 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__2867  (.I0(\edb_top_inst/n1852 ), .I1(\edb_top_inst/edb_user_dr[32] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2867 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2868  (.I0(\edb_top_inst/edb_user_dr[33] ), 
            .I1(\edb_top_inst/la0/word_count[4] ), .I2(\edb_top_inst/n1796 ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2868 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__2869  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/n1796 ), .O(\edb_top_inst/n1853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2869 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2870  (.I0(\edb_top_inst/edb_user_dr[34] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/n1853 ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2870 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__2871  (.I0(\edb_top_inst/la0/word_count[5] ), 
            .I1(\edb_top_inst/n1853 ), .O(\edb_top_inst/n1854 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2871 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2872  (.I0(\edb_top_inst/edb_user_dr[35] ), 
            .I1(\edb_top_inst/la0/word_count[6] ), .I2(\edb_top_inst/n1854 ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2872 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__2873  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/la0/word_count[6] ), 
            .I3(\edb_top_inst/n1796 ), .O(\edb_top_inst/n1855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2873 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__2874  (.I0(\edb_top_inst/edb_user_dr[36] ), 
            .I1(\edb_top_inst/la0/word_count[7] ), .I2(\edb_top_inst/n1855 ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2874 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__2875  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/n1855 ), .O(\edb_top_inst/n1856 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2875 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2876  (.I0(\edb_top_inst/edb_user_dr[37] ), 
            .I1(\edb_top_inst/la0/word_count[8] ), .I2(\edb_top_inst/n1856 ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2876 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__2877  (.I0(\edb_top_inst/la0/word_count[8] ), 
            .I1(\edb_top_inst/n1856 ), .O(\edb_top_inst/n1857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2877 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2878  (.I0(\edb_top_inst/edb_user_dr[38] ), 
            .I1(\edb_top_inst/la0/word_count[9] ), .I2(\edb_top_inst/n1857 ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2878 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__2879  (.I0(\edb_top_inst/la0/word_count[7] ), 
            .I1(\edb_top_inst/la0/word_count[8] ), .I2(\edb_top_inst/la0/word_count[9] ), 
            .I3(\edb_top_inst/n1855 ), .O(\edb_top_inst/n1858 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2879 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__2880  (.I0(\edb_top_inst/edb_user_dr[39] ), 
            .I1(\edb_top_inst/la0/word_count[10] ), .I2(\edb_top_inst/n1858 ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2880 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__2881  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/n1858 ), .I2(\edb_top_inst/la0/word_count[11] ), 
            .O(\edb_top_inst/n1859 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2881 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__2882  (.I0(\edb_top_inst/n1859 ), .I1(\edb_top_inst/edb_user_dr[40] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2882 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2883  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/la0/word_count[11] ), .I2(\edb_top_inst/n1858 ), 
            .O(\edb_top_inst/n1860 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2883 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__2884  (.I0(\edb_top_inst/edb_user_dr[41] ), 
            .I1(\edb_top_inst/la0/word_count[12] ), .I2(\edb_top_inst/n1860 ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2884 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__2885  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/n1860 ), .I2(\edb_top_inst/la0/word_count[13] ), 
            .O(\edb_top_inst/n1861 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2885 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__2886  (.I0(\edb_top_inst/n1861 ), .I1(\edb_top_inst/edb_user_dr[42] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2886 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2887  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/la0/word_count[13] ), .I2(\edb_top_inst/n1860 ), 
            .O(\edb_top_inst/n1862 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2887 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__2888  (.I0(\edb_top_inst/edb_user_dr[43] ), 
            .I1(\edb_top_inst/la0/word_count[14] ), .I2(\edb_top_inst/n1862 ), 
            .I3(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2888 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__2889  (.I0(\edb_top_inst/la0/word_count[14] ), 
            .I1(\edb_top_inst/n1862 ), .I2(\edb_top_inst/la0/word_count[15] ), 
            .O(\edb_top_inst/n1863 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2889 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__2890  (.I0(\edb_top_inst/n1863 ), .I1(\edb_top_inst/edb_user_dr[44] ), 
            .I2(\edb_top_inst/n1768 ), .O(\edb_top_inst/la0/data_to_word_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2890 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__2891  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/n1827 ), 
            .O(\edb_top_inst/n1864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2891 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__2892  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[1] ), .I2(\edb_top_inst/n1864 ), 
            .O(\edb_top_inst/n1865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2892 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__2893  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n1866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb8f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2893 .LUTMASK = 16'hfb8f;
    EFX_LUT4 \edb_top_inst/LUT__2894  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n1826 ), .O(\edb_top_inst/n1867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2894 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2895  (.I0(\edb_top_inst/n1867 ), .I1(\edb_top_inst/la0/internal_register_select[3] ), 
            .I2(\edb_top_inst/n1802 ), .O(\edb_top_inst/n1868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2895 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__2896  (.I0(\edb_top_inst/n1866 ), .I1(\edb_top_inst/la0/data_from_biu[1] ), 
            .I2(\edb_top_inst/n1868 ), .I3(\edb_top_inst/n1802 ), .O(\edb_top_inst/n1869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2896 .LUTMASK = 16'h0c05;
    EFX_LUT4 \edb_top_inst/LUT__2897  (.I0(\edb_top_inst/n1869 ), .I1(\edb_top_inst/n1865 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[2] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2897 .LUTMASK = 16'heef0;
    EFX_LUT4 \edb_top_inst/LUT__2898  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/n1826 ), 
            .O(\edb_top_inst/n1870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2898 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__2899  (.I0(\edb_top_inst/n1870 ), .I1(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I2(\edb_top_inst/n1867 ), .I3(\edb_top_inst/n1802 ), .O(\edb_top_inst/n1871 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2899 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__2900  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n1872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2900 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2901  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/n1872 ), 
            .O(\edb_top_inst/n1873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2901 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__2902  (.I0(\edb_top_inst/n1873 ), .I1(\edb_top_inst/la0/data_from_biu[2] ), 
            .I2(\edb_top_inst/n1868 ), .I3(\edb_top_inst/n1802 ), .O(\edb_top_inst/n1874 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2902 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__2903  (.I0(\edb_top_inst/n1874 ), .I1(\edb_top_inst/n1871 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[3] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2903 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__2904  (.I0(\edb_top_inst/n1826 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .I2(\edb_top_inst/la0/internal_register_select[3] ), .I3(\edb_top_inst/n1802 ), 
            .O(\edb_top_inst/n1875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2904 .LUTMASK = 16'h007d;
    EFX_LUT4 \edb_top_inst/LUT__2905  (.I0(\edb_top_inst/n1875 ), .I1(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/n1876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2905 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2906  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n1802 ), .I2(\edb_top_inst/n1756 ), .I3(\edb_top_inst/n1814 ), 
            .O(\edb_top_inst/n1877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2906 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__2907  (.I0(\edb_top_inst/la0/la_trig_mask[3] ), 
            .I1(\edb_top_inst/n1870 ), .I2(\edb_top_inst/la0/data_out_shift_reg[4] ), 
            .I3(\edb_top_inst/n1877 ), .O(\edb_top_inst/n1878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2907 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__2908  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(\edb_top_inst/la0/data_from_biu[3] ), .I2(\edb_top_inst/n1877 ), 
            .O(\edb_top_inst/n1879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2908 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2909  (.I0(\edb_top_inst/n1868 ), .I1(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/n1880 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2909 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2910  (.I0(\edb_top_inst/n1879 ), .I1(\edb_top_inst/n1880 ), 
            .I2(\edb_top_inst/n1876 ), .I3(\edb_top_inst/n1878 ), .O(\edb_top_inst/la0/n2440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2910 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__2911  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/data_from_biu[4] ), .I2(\edb_top_inst/n1802 ), 
            .O(\edb_top_inst/n1881 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2911 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2912  (.I0(\edb_top_inst/la0/la_trig_mask[4] ), 
            .I1(\edb_top_inst/n1870 ), .I2(\edb_top_inst/la0/data_out_shift_reg[5] ), 
            .I3(\edb_top_inst/n1877 ), .O(\edb_top_inst/n1882 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2912 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__2913  (.I0(\edb_top_inst/n1882 ), .I1(\edb_top_inst/n1881 ), 
            .I2(\edb_top_inst/n1880 ), .O(\edb_top_inst/la0/n2439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2913 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2914  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(\edb_top_inst/la0/data_from_biu[5] ), .I2(\edb_top_inst/n1802 ), 
            .O(\edb_top_inst/n1883 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2914 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2915  (.I0(\edb_top_inst/la0/la_trig_mask[5] ), 
            .I1(\edb_top_inst/n1870 ), .I2(\edb_top_inst/la0/data_out_shift_reg[6] ), 
            .I3(\edb_top_inst/n1877 ), .O(\edb_top_inst/n1884 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2915 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__2916  (.I0(\edb_top_inst/n1884 ), .I1(\edb_top_inst/n1883 ), 
            .I2(\edb_top_inst/n1880 ), .O(\edb_top_inst/la0/n2438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2916 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2917  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[6] ), .I2(\edb_top_inst/n1864 ), 
            .O(\edb_top_inst/n1885 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2917 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__2918  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(\edb_top_inst/la0/data_from_biu[6] ), .I2(\edb_top_inst/n1877 ), 
            .I3(\edb_top_inst/n1880 ), .O(\edb_top_inst/n1886 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2918 .LUTMASK = 16'hac00;
    EFX_LUT4 \edb_top_inst/LUT__2919  (.I0(\edb_top_inst/n1885 ), .I1(\edb_top_inst/la0/data_out_shift_reg[7] ), 
            .I2(\edb_top_inst/n1886 ), .I3(\edb_top_inst/n1831 ), .O(\edb_top_inst/la0/n2437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfafc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2919 .LUTMASK = 16'hfafc;
    EFX_LUT4 \edb_top_inst/LUT__2920  (.I0(\edb_top_inst/la0/la_trig_mask[7] ), 
            .I1(\edb_top_inst/n1870 ), .I2(\edb_top_inst/la0/data_out_shift_reg[8] ), 
            .I3(\edb_top_inst/n1877 ), .O(\edb_top_inst/n1887 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2920 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__2921  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(\edb_top_inst/la0/data_from_biu[7] ), .I2(\edb_top_inst/n1877 ), 
            .O(\edb_top_inst/n1888 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2921 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2922  (.I0(\edb_top_inst/n1888 ), .I1(\edb_top_inst/n1880 ), 
            .I2(\edb_top_inst/n1876 ), .I3(\edb_top_inst/n1887 ), .O(\edb_top_inst/la0/n2436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2922 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__2923  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(\edb_top_inst/la0/data_from_biu[8] ), .I2(\edb_top_inst/n1802 ), 
            .O(\edb_top_inst/n1889 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2923 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2924  (.I0(\edb_top_inst/la0/la_trig_mask[8] ), 
            .I1(\edb_top_inst/n1870 ), .I2(\edb_top_inst/la0/data_out_shift_reg[9] ), 
            .I3(\edb_top_inst/n1877 ), .O(\edb_top_inst/n1890 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2924 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__2925  (.I0(\edb_top_inst/n1890 ), .I1(\edb_top_inst/n1889 ), 
            .I2(\edb_top_inst/n1880 ), .O(\edb_top_inst/la0/n2435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2925 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2926  (.I0(\edb_top_inst/n1870 ), .I1(\edb_top_inst/la0/la_trig_mask[9] ), 
            .I2(\edb_top_inst/n1867 ), .I3(\edb_top_inst/n1802 ), .O(\edb_top_inst/n1891 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2926 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__2927  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(\edb_top_inst/la0/data_from_biu[9] ), .I2(\edb_top_inst/n1868 ), 
            .I3(\edb_top_inst/n1802 ), .O(\edb_top_inst/n1892 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2927 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__2928  (.I0(\edb_top_inst/n1892 ), .I1(\edb_top_inst/n1891 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[10] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h11f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2928 .LUTMASK = 16'h11f0;
    EFX_LUT4 \edb_top_inst/LUT__2929  (.I0(\edb_top_inst/la0/la_trig_mask[10] ), 
            .I1(\edb_top_inst/n1870 ), .I2(\edb_top_inst/la0/data_out_shift_reg[11] ), 
            .I3(\edb_top_inst/n1877 ), .O(\edb_top_inst/n1893 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2929 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__2930  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(\edb_top_inst/la0/data_from_biu[10] ), .I2(\edb_top_inst/n1877 ), 
            .O(\edb_top_inst/n1894 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2930 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2931  (.I0(\edb_top_inst/n1894 ), .I1(\edb_top_inst/n1880 ), 
            .I2(\edb_top_inst/n1876 ), .I3(\edb_top_inst/n1893 ), .O(\edb_top_inst/la0/n2433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2931 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__2932  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[11] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1895 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2932 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__2933  (.I0(\edb_top_inst/n1895 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[12] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2933 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2934  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[12] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1896 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2934 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2935  (.I0(\edb_top_inst/n1896 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[13] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2935 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2936  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[13] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1897 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2936 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2937  (.I0(\edb_top_inst/n1897 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[14] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2937 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2938  (.I0(\edb_top_inst/la0/la_sample_cnt[11] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[14] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1898 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2938 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__2939  (.I0(\edb_top_inst/n1898 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[15] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2939 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2940  (.I0(\edb_top_inst/la0/la_sample_cnt[12] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[15] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1899 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2940 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2941  (.I0(\edb_top_inst/n1899 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[16] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2941 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2942  (.I0(\edb_top_inst/la0/la_trig_mask[16] ), 
            .I1(\edb_top_inst/n1870 ), .O(\edb_top_inst/n1900 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2942 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__2943  (.I0(\edb_top_inst/n1900 ), .I1(\edb_top_inst/n1864 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[17] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2943 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2944  (.I0(\edb_top_inst/la0/la_trig_mask[17] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n1901 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2944 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2945  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n1827 ), .O(\edb_top_inst/n1902 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2945 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__2946  (.I0(\edb_top_inst/n1901 ), .I1(\edb_top_inst/n1902 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[18] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2946 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2947  (.I0(\edb_top_inst/la0/la_trig_mask[18] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n1903 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2947 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__2948  (.I0(\edb_top_inst/n1903 ), .I1(\edb_top_inst/n1902 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[19] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2948 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2949  (.I0(\edb_top_inst/n1870 ), .I1(\edb_top_inst/la0/la_trig_mask[19] ), 
            .I2(\edb_top_inst/n1867 ), .O(\edb_top_inst/n1904 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2949 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__2950  (.I0(\edb_top_inst/n1904 ), .I1(\edb_top_inst/n1868 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[20] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2950 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2951  (.I0(\edb_top_inst/la0/la_trig_mask[20] ), 
            .I1(\edb_top_inst/la0/la_run_trig ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1905 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2951 .LUTMASK = 16'h05f3;
    EFX_LUT4 \edb_top_inst/LUT__2952  (.I0(\edb_top_inst/n1905 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[21] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2952 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2953  (.I0(\edb_top_inst/la0/la_trig_mask[21] ), 
            .I1(\edb_top_inst/la0/la_run_trig_imdt ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1906 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2953 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2954  (.I0(\edb_top_inst/n1906 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[22] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2954 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2955  (.I0(\edb_top_inst/la0/la_trig_mask[22] ), 
            .I1(\edb_top_inst/la0/la_stop_trig ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1907 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2955 .LUTMASK = 16'h0503;
    EFX_LUT4 \edb_top_inst/LUT__2956  (.I0(\edb_top_inst/n1907 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[23] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2956 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2957  (.I0(\edb_top_inst/la0/la_trig_mask[23] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[0] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1908 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2957 .LUTMASK = 16'h05f3;
    EFX_LUT4 \edb_top_inst/LUT__2958  (.I0(\edb_top_inst/n1908 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[24] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2958 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2959  (.I0(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[24] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1909 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2959 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__2960  (.I0(\edb_top_inst/n1909 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[25] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2960 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2961  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[25] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1910 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2961 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2962  (.I0(\edb_top_inst/n1910 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[26] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2962 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2963  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[26] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1911 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2963 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__2964  (.I0(\edb_top_inst/n1911 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[27] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2964 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2965  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[27] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1912 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2965 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2966  (.I0(\edb_top_inst/n1912 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[28] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2966 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2967  (.I0(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[28] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1913 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2967 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2968  (.I0(\edb_top_inst/n1913 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[29] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2968 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2969  (.I0(\edb_top_inst/la0/la_trig_mask[29] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[6] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1914 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2969 .LUTMASK = 16'h05f3;
    EFX_LUT4 \edb_top_inst/LUT__2970  (.I0(\edb_top_inst/n1914 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[30] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2970 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2971  (.I0(\edb_top_inst/la0/la_trig_mask[30] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[7] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1915 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2971 .LUTMASK = 16'h05f3;
    EFX_LUT4 \edb_top_inst/LUT__2972  (.I0(\edb_top_inst/n1915 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[31] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2972 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2973  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[31] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1916 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2973 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2974  (.I0(\edb_top_inst/n1916 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[32] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2974 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2975  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[32] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1917 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2975 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__2976  (.I0(\edb_top_inst/n1917 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[33] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2976 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2977  (.I0(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[33] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1918 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2977 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2978  (.I0(\edb_top_inst/n1918 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[34] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2978 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2979  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[34] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1919 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2979 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2980  (.I0(\edb_top_inst/n1919 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[35] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2980 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2981  (.I0(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[35] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1920 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2981 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__2982  (.I0(\edb_top_inst/n1920 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[36] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2982 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2983  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[36] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1921 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2983 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__2984  (.I0(\edb_top_inst/n1921 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[37] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2984 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2985  (.I0(\edb_top_inst/la0/la_trig_mask[37] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[14] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1922 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2985 .LUTMASK = 16'h05f3;
    EFX_LUT4 \edb_top_inst/LUT__2986  (.I0(\edb_top_inst/n1922 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[38] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2986 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2987  (.I0(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[38] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1923 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2987 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__2988  (.I0(\edb_top_inst/n1923 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[39] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2988 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2989  (.I0(\edb_top_inst/la0/la_trig_mask[39] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[16] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1924 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2989 .LUTMASK = 16'h05f3;
    EFX_LUT4 \edb_top_inst/LUT__2990  (.I0(\edb_top_inst/n1924 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[40] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2990 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2991  (.I0(\edb_top_inst/la0/la_trig_mask[40] ), 
            .I1(\edb_top_inst/la0/la_trig_pattern[0] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1925 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2991 .LUTMASK = 16'h05f3;
    EFX_LUT4 \edb_top_inst/LUT__2992  (.I0(\edb_top_inst/n1925 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[41] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2992 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2993  (.I0(\edb_top_inst/la0/la_trig_mask[41] ), 
            .I1(\edb_top_inst/la0/la_trig_pattern[1] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n1926 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2993 .LUTMASK = 16'h05f3;
    EFX_LUT4 \edb_top_inst/LUT__2994  (.I0(\edb_top_inst/n1926 ), .I1(\edb_top_inst/n1827 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[42] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2994 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2995  (.I0(\edb_top_inst/la0/la_trig_mask[42] ), 
            .I1(\edb_top_inst/la0/la_capture_pattern[0] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1927 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2995 .LUTMASK = 16'h5353;
    EFX_LUT4 \edb_top_inst/LUT__2996  (.I0(\edb_top_inst/n1927 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[43] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2401 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2996 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2997  (.I0(\edb_top_inst/la0/la_capture_pattern[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[43] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n1928 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2997 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__2998  (.I0(\edb_top_inst/n1928 ), .I1(\edb_top_inst/n1828 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[44] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2998 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__2999  (.I0(\edb_top_inst/n1870 ), .I1(\edb_top_inst/n1877 ), 
            .O(\edb_top_inst/n1929 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2999 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3000  (.I0(\edb_top_inst/n1831 ), .I1(\edb_top_inst/la0/data_out_shift_reg[45] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[44] ), .I3(\edb_top_inst/n1929 ), 
            .O(\edb_top_inst/la0/n2399 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3000 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3001  (.I0(\edb_top_inst/n1831 ), .I1(\edb_top_inst/la0/data_out_shift_reg[46] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[45] ), .I3(\edb_top_inst/n1929 ), 
            .O(\edb_top_inst/la0/n2398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3001 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3002  (.I0(\edb_top_inst/n1831 ), .I1(\edb_top_inst/la0/data_out_shift_reg[47] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[46] ), .I3(\edb_top_inst/n1929 ), 
            .O(\edb_top_inst/la0/n2397 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3002 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3003  (.I0(\edb_top_inst/n1870 ), .I1(\edb_top_inst/la0/la_trig_mask[47] ), 
            .I2(\edb_top_inst/n1867 ), .O(\edb_top_inst/n1930 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3003 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3004  (.I0(\edb_top_inst/n1930 ), .I1(\edb_top_inst/n1868 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[48] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3004 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3005  (.I0(\edb_top_inst/n1831 ), .I1(\edb_top_inst/la0/data_out_shift_reg[49] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[48] ), .I3(\edb_top_inst/n1929 ), 
            .O(\edb_top_inst/la0/n2395 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3005 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3006  (.I0(\edb_top_inst/n1831 ), .I1(\edb_top_inst/la0/data_out_shift_reg[50] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[49] ), .I3(\edb_top_inst/n1929 ), 
            .O(\edb_top_inst/la0/n2394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3006 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3007  (.I0(\edb_top_inst/n1870 ), .I1(\edb_top_inst/la0/la_trig_mask[50] ), 
            .I2(\edb_top_inst/n1867 ), .O(\edb_top_inst/n1931 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3007 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3008  (.I0(\edb_top_inst/n1931 ), .I1(\edb_top_inst/n1868 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[51] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2393 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3008 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3009  (.I0(\edb_top_inst/la0/la_trig_mask[51] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n1932 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3009 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3010  (.I0(\edb_top_inst/n1932 ), .I1(\edb_top_inst/n1902 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[52] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3010 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3011  (.I0(\edb_top_inst/la0/la_trig_mask[52] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n1933 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3011 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3012  (.I0(\edb_top_inst/n1933 ), .I1(\edb_top_inst/n1902 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[53] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2391 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3012 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3013  (.I0(\edb_top_inst/la0/la_trig_mask[53] ), 
            .I1(\edb_top_inst/n1870 ), .O(\edb_top_inst/n1934 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3013 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3014  (.I0(\edb_top_inst/n1934 ), .I1(\edb_top_inst/n1864 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[54] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3014 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3015  (.I0(\edb_top_inst/la0/la_trig_mask[54] ), 
            .I1(\edb_top_inst/n1870 ), .O(\edb_top_inst/n1935 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3015 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3016  (.I0(\edb_top_inst/n1935 ), .I1(\edb_top_inst/n1864 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[55] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2389 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3016 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3017  (.I0(\edb_top_inst/la0/la_trig_mask[55] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n1936 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3017 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3018  (.I0(\edb_top_inst/n1936 ), .I1(\edb_top_inst/n1902 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[56] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2388 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3018 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3019  (.I0(\edb_top_inst/la0/la_trig_mask[56] ), 
            .I1(\edb_top_inst/n1870 ), .O(\edb_top_inst/n1937 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3019 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3020  (.I0(\edb_top_inst/n1937 ), .I1(\edb_top_inst/n1864 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[57] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2387 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3020 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3021  (.I0(\edb_top_inst/n1831 ), .I1(\edb_top_inst/la0/data_out_shift_reg[58] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[57] ), .I3(\edb_top_inst/n1929 ), 
            .O(\edb_top_inst/la0/n2386 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3021 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3022  (.I0(\edb_top_inst/n1870 ), .I1(\edb_top_inst/la0/la_trig_mask[58] ), 
            .I2(\edb_top_inst/n1867 ), .O(\edb_top_inst/n1938 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3022 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3023  (.I0(\edb_top_inst/n1938 ), .I1(\edb_top_inst/n1868 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[59] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2385 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3023 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3024  (.I0(\edb_top_inst/la0/la_trig_mask[59] ), 
            .I1(\edb_top_inst/n1870 ), .O(\edb_top_inst/n1939 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3024 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3025  (.I0(\edb_top_inst/n1939 ), .I1(\edb_top_inst/n1864 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[60] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2384 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3025 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3026  (.I0(\edb_top_inst/la0/la_trig_mask[60] ), 
            .I1(\edb_top_inst/n1870 ), .O(\edb_top_inst/n1940 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3026 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3027  (.I0(\edb_top_inst/n1940 ), .I1(\edb_top_inst/n1864 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[61] ), .I3(\edb_top_inst/n1831 ), 
            .O(\edb_top_inst/la0/n2383 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3027 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3028  (.I0(\edb_top_inst/n1831 ), .I1(\edb_top_inst/la0/data_out_shift_reg[62] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[61] ), .I3(\edb_top_inst/n1929 ), 
            .O(\edb_top_inst/la0/n2382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3028 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3029  (.I0(\edb_top_inst/n1831 ), .I1(\edb_top_inst/la0/data_out_shift_reg[63] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[62] ), .I3(\edb_top_inst/n1929 ), 
            .O(\edb_top_inst/la0/n2381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3029 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3030  (.I0(\edb_top_inst/n1870 ), .I1(\edb_top_inst/la0/la_trig_mask[63] ), 
            .I2(\edb_top_inst/n1867 ), .O(\edb_top_inst/n1941 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3030 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3031  (.I0(\edb_top_inst/n1941 ), .I1(\edb_top_inst/n1868 ), 
            .I2(\edb_top_inst/n1831 ), .O(\edb_top_inst/la0/n2380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3031 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3032  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/n1761 ), .O(\edb_top_inst/n1942 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3032 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3033  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .I2(\edb_top_inst/n1817 ), 
            .I3(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n1943 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3033 .LUTMASK = 16'hf100;
    EFX_LUT4 \edb_top_inst/LUT__3034  (.I0(\edb_top_inst/n1814 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/n1798 ), .I3(\edb_top_inst/n1943 ), .O(\edb_top_inst/n1944 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3034 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__3035  (.I0(\edb_top_inst/n1944 ), .I1(\edb_top_inst/n1942 ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/la0/module_next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3035 .LUTMASK = 16'hc5c5;
    EFX_LUT4 \edb_top_inst/LUT__3036  (.I0(\edb_top_inst/n1756 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n1945 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3036 .LUTMASK = 16'hd3d3;
    EFX_LUT4 \edb_top_inst/LUT__3037  (.I0(\edb_top_inst/n1818 ), .I1(\edb_top_inst/n1795 ), 
            .I2(\edb_top_inst/n1797 ), .I3(\edb_top_inst/n1945 ), .O(\edb_top_inst/n1946 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7770, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3037 .LUTMASK = 16'h7770;
    EFX_LUT4 \edb_top_inst/LUT__3038  (.I0(\edb_top_inst/n1804 ), .I1(\edb_top_inst/n1946 ), 
            .I2(jtag_inst1_UPDATE), .I3(\edb_top_inst/n1761 ), .O(\edb_top_inst/la0/module_next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h330b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3038 .LUTMASK = 16'h330b;
    EFX_LUT4 \edb_top_inst/LUT__3039  (.I0(\edb_top_inst/n1788 ), .I1(\edb_top_inst/n1811 ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n1947 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf70f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3039 .LUTMASK = 16'hf70f;
    EFX_LUT4 \edb_top_inst/LUT__3040  (.I0(\edb_top_inst/n1797 ), .I1(\edb_top_inst/n1756 ), 
            .I2(jtag_inst1_UPDATE), .I3(\edb_top_inst/n1947 ), .O(\edb_top_inst/la0/module_next_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3040 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__3041  (.I0(\edb_top_inst/la0/crc_data_out[1] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3041 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3042  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/n1761 ), .I2(\edb_top_inst/la0/module_state[3] ), 
            .I3(\edb_top_inst/n1810 ), .O(\edb_top_inst/ceg_net221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3042 .LUTMASK = 16'hbf00;
    EFX_LUT4 \edb_top_inst/LUT__3043  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3043 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3044  (.I0(\edb_top_inst/la0/crc_data_out[3] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3044 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3045  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3045 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3046  (.I0(\edb_top_inst/la0/crc_data_out[5] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3046 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3047  (.I0(jtag_inst1_TDI), .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/crc_data_out[0] ), 
            .O(\edb_top_inst/n1948 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3047 .LUTMASK = 16'hac53;
    EFX_LUT4 \edb_top_inst/LUT__3048  (.I0(\edb_top_inst/n1948 ), .I1(\edb_top_inst/n1809 ), 
            .O(\edb_top_inst/n1949 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3048 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3049  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[6] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3049 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3051  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3051 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__2677  (.I0(\edb_top_inst/la0/crc_data_out[10] ), 
            .I1(\edb_top_inst/edb_user_dr[60] ), .I2(\edb_top_inst/la0/crc_data_out[11] ), 
            .I3(\edb_top_inst/edb_user_dr[61] ), .O(\edb_top_inst/n1730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__2677 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3052  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3052 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3053  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[9] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3053 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3054  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[10] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3054 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3055  (.I0(\edb_top_inst/la0/crc_data_out[11] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3055 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3056  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3056 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3057  (.I0(\edb_top_inst/la0/crc_data_out[13] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3057 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3058  (.I0(\edb_top_inst/la0/crc_data_out[14] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3058 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3059  (.I0(\edb_top_inst/la0/crc_data_out[15] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3059 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3060  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[16] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3060 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3061  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3061 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3062  (.I0(\edb_top_inst/la0/crc_data_out[18] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3062 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3063  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3063 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3064  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[20] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3064 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3065  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[21] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3065 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3066  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[22] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3066 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3067  (.I0(\edb_top_inst/la0/crc_data_out[23] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3067 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3068  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[24] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3068 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3069  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[25] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3069 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3070  (.I0(\edb_top_inst/la0/crc_data_out[26] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3070 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3071  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[27] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3071 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3072  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[28] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3072 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3073  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/n1780 ), .O(\edb_top_inst/la0/axi_crc_i/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3073 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3074  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[30] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3074 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3075  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[31] ), .I2(\edb_top_inst/n1949 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3075 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3076  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n1949 ), .O(\edb_top_inst/la0/axi_crc_i/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3076 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3077  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3077 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3078  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3078 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3079  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n16 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n17 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3079 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3080  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3080 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__3081  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n1950 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3081 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__3082  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n1950 ), .O(\edb_top_inst/n1951 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3082 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__3083  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n1952 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3083 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__3084  (.I0(\edb_top_inst/n1952 ), .I1(\edb_top_inst/n1951 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3084 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3085  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3085 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3086  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3086 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3087  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n16 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n17 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3087 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3088  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3088 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__3089  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n1953 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3089 .LUTMASK = 16'h503f;
    EFX_LUT4 \edb_top_inst/LUT__3090  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n1953 ), .O(\edb_top_inst/n1954 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3090 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__3091  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n1955 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3091 .LUTMASK = 16'h035f;
    EFX_LUT4 \edb_top_inst/LUT__3092  (.I0(\edb_top_inst/n1955 ), .I1(\edb_top_inst/n1954 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3092 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3093  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3093 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3094  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3094 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3095  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), .O(\edb_top_inst/n1956 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3095 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3096  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n1957 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3096 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3097  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), 
            .I1(\edb_top_inst/n1956 ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n1957 ), .O(\edb_top_inst/n1958 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3097 .LUTMASK = 16'h7100;
    EFX_LUT4 \edb_top_inst/LUT__3098  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/n1959 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3098 .LUTMASK = 16'h8eaf;
    EFX_LUT4 \edb_top_inst/LUT__3099  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/n1958 ), .I3(\edb_top_inst/n1959 ), .O(\edb_top_inst/n1960 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3099 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__3100  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/n1960 ), .O(\edb_top_inst/n1961 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3100 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__3101  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/n1961 ), .O(\edb_top_inst/n1962 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3101 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__3102  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I2(\edb_top_inst/n1962 ), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3102 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__3103  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n1963 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3103 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3104  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/n1964 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3104 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3105  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n1965 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3105 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3106  (.I0(\edb_top_inst/n1957 ), .I1(\edb_top_inst/n1963 ), 
            .I2(\edb_top_inst/n1964 ), .I3(\edb_top_inst/n1965 ), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3106 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__3107  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n1966 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3107 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__3108  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n1967 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3108 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3109  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n1968 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3109 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3110  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n1969 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3110 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3111  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n1970 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3111 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3112  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n1971 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3112 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3113  (.I0(\edb_top_inst/n1968 ), .I1(\edb_top_inst/n1969 ), 
            .I2(\edb_top_inst/n1970 ), .I3(\edb_top_inst/n1971 ), .O(\edb_top_inst/n1972 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3113 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3114  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/n1967 ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n1972 ), .O(\edb_top_inst/n1973 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h752f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3114 .LUTMASK = 16'h752f;
    EFX_LUT4 \edb_top_inst/LUT__3115  (.I0(\edb_top_inst/n1973 ), .I1(\edb_top_inst/n1966 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3115 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3116  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3116 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3117  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3117 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3118  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3118 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3119  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3119 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3120  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3120 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3121  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3121 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3122  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3122 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3123  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3123 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3124  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3124 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3125  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3125 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3126  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3126 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3127  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3127 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3128  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3128 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3129  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3129 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3130  (.I0(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n1974 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3130 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3131  (.I0(\edb_top_inst/n1974 ), .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[0] ), .I3(\edb_top_inst/la0/la_trig_pattern[0] ), 
            .O(\edb_top_inst/n1975 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2acf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3131 .LUTMASK = 16'h2acf;
    EFX_LUT4 \edb_top_inst/LUT__3132  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[2] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[1] ), .O(\edb_top_inst/n1976 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3132 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__3133  (.I0(\edb_top_inst/n1976 ), .I1(\edb_top_inst/la0/la_trig_pattern[0] ), 
            .I2(\edb_top_inst/la0/la_trig_pattern[1] ), .I3(\edb_top_inst/n1975 ), 
            .O(\edb_top_inst/n1977 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2dc3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3133 .LUTMASK = 16'h2dc3;
    EFX_LUT4 \edb_top_inst/LUT__3134  (.I0(\edb_top_inst/la0/la_trig_mask[0] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[1] ), .I2(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I3(\edb_top_inst/n1977 ), .O(\edb_top_inst/la0/trigger_tu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3134 .LUTMASK = 16'h00fe;
    EFX_LUT4 \edb_top_inst/LUT__3135  (.I0(\edb_top_inst/la0/tu_trigger ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n1978 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3135 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3136  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n1979 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3136 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3137  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(\edb_top_inst/n1979 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .O(\edb_top_inst/n1980 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3137 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__3138  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n1981 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3138 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3139  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n1982 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3139 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3140  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), .I2(\edb_top_inst/n1982 ), 
            .I3(\edb_top_inst/n1981 ), .O(\edb_top_inst/n1983 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3140 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__3141  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n1984 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3141 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__3142  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(\edb_top_inst/n1984 ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I3(\edb_top_inst/n1983 ), .O(\edb_top_inst/n1985 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3142 .LUTMASK = 16'he100;
    EFX_LUT4 \edb_top_inst/LUT__3143  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n1986 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3143 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3144  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n1987 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3144 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3145  (.I0(\edb_top_inst/n1986 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I3(\edb_top_inst/n1987 ), 
            .O(\edb_top_inst/n1988 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3145 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__3146  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n1989 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3146 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__3147  (.I0(\edb_top_inst/n1989 ), .I1(\edb_top_inst/n1981 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), .O(\edb_top_inst/n1990 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3147 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__3148  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n1984 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] ), 
            .O(\edb_top_inst/n1991 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf807, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3148 .LUTMASK = 16'hf807;
    EFX_LUT4 \edb_top_inst/LUT__3149  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n1992 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3149 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3150  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n1992 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), .O(\edb_top_inst/n1993 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf20d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3150 .LUTMASK = 16'hf20d;
    EFX_LUT4 \edb_top_inst/LUT__3151  (.I0(\edb_top_inst/n1988 ), .I1(\edb_top_inst/n1990 ), 
            .I2(\edb_top_inst/n1991 ), .I3(\edb_top_inst/n1993 ), .O(\edb_top_inst/n1994 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3151 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3152  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n1995 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3152 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3153  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n1996 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3153 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3154  (.I0(\edb_top_inst/n1995 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .I3(\edb_top_inst/n1996 ), 
            .O(\edb_top_inst/n1997 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3154 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__3155  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n1998 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3155 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3156  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n1999 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3156 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3157  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n1998 ), .I2(\edb_top_inst/n1999 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .O(\edb_top_inst/n2000 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3157 .LUTMASK = 16'h40bf;
    EFX_LUT4 \edb_top_inst/LUT__3158  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n2001 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3158 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__3159  (.I0(\edb_top_inst/n1997 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I2(\edb_top_inst/n2000 ), .I3(\edb_top_inst/n2001 ), .O(\edb_top_inst/n2002 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1004, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3159 .LUTMASK = 16'h1004;
    EFX_LUT4 \edb_top_inst/LUT__3160  (.I0(\edb_top_inst/n1980 ), .I1(\edb_top_inst/n1985 ), 
            .I2(\edb_top_inst/n1994 ), .I3(\edb_top_inst/n2002 ), .O(\edb_top_inst/n2003 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3160 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3161  (.I0(\edb_top_inst/n2003 ), .I1(\edb_top_inst/n1978 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n2004 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3161 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3162  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n2005 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3162 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3163  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/n2004 ), .I2(\edb_top_inst/n2005 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n2006 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3163 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__3164  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n1986 ), .I2(\edb_top_inst/n1981 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .O(\edb_top_inst/n2007 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h807f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3164 .LUTMASK = 16'h807f;
    EFX_LUT4 \edb_top_inst/LUT__3165  (.I0(\edb_top_inst/n1992 ), .I1(\edb_top_inst/n1981 ), 
            .I2(\edb_top_inst/n2007 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .O(\edb_top_inst/n2008 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b04, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3165 .LUTMASK = 16'h0b04;
    EFX_LUT4 \edb_top_inst/LUT__3166  (.I0(\edb_top_inst/n1996 ), .I1(\edb_top_inst/n1998 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .O(\edb_top_inst/n2009 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3166 .LUTMASK = 16'h8f70;
    EFX_LUT4 \edb_top_inst/LUT__3167  (.I0(\edb_top_inst/n1990 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I2(\edb_top_inst/n2009 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .O(\edb_top_inst/n2010 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3167 .LUTMASK = 16'h0c05;
    EFX_LUT4 \edb_top_inst/LUT__3168  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n2011 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3168 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3169  (.I0(\edb_top_inst/n2011 ), .I1(\edb_top_inst/n1995 ), 
            .I2(\edb_top_inst/n2001 ), .O(\edb_top_inst/n2012 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3169 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3170  (.I0(\edb_top_inst/n1993 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), .I3(\edb_top_inst/n2012 ), 
            .O(\edb_top_inst/n2013 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3170 .LUTMASK = 16'hf53f;
    EFX_LUT4 \edb_top_inst/LUT__3171  (.I0(\edb_top_inst/n2013 ), .I1(\edb_top_inst/n2010 ), 
            .I2(\edb_top_inst/n2008 ), .O(\edb_top_inst/n2014 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3171 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3172  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n1984 ), .O(\edb_top_inst/n2015 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3172 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3173  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n2016 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1ffe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3173 .LUTMASK = 16'h1ffe;
    EFX_LUT4 \edb_top_inst/LUT__3174  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n2016 ), .O(\edb_top_inst/n2017 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3174 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3175  (.I0(\edb_top_inst/n2015 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), .I3(\edb_top_inst/n2017 ), 
            .O(\edb_top_inst/n2018 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3175 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__3176  (.I0(\edb_top_inst/n1995 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), .I3(\edb_top_inst/n1996 ), 
            .O(\edb_top_inst/n2019 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ecf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3176 .LUTMASK = 16'h7ecf;
    EFX_LUT4 \edb_top_inst/LUT__3177  (.I0(\edb_top_inst/n1992 ), .I1(\edb_top_inst/n1979 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n2020 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3177 .LUTMASK = 16'h0c05;
    EFX_LUT4 \edb_top_inst/LUT__3178  (.I0(\edb_top_inst/n1987 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), .I3(\edb_top_inst/n2020 ), 
            .O(\edb_top_inst/n2021 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3178 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__3179  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n1992 ), .I2(\edb_top_inst/n1982 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .O(\edb_top_inst/n2022 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3179 .LUTMASK = 16'hb04f;
    EFX_LUT4 \edb_top_inst/LUT__3180  (.I0(\edb_top_inst/n2018 ), .I1(\edb_top_inst/n2019 ), 
            .I2(\edb_top_inst/n2021 ), .I3(\edb_top_inst/n2022 ), .O(\edb_top_inst/n2023 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3180 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3181  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/n1982 ), 
            .O(\edb_top_inst/n2024 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3181 .LUTMASK = 16'h0e0e;
    EFX_LUT4 \edb_top_inst/LUT__3182  (.I0(\edb_top_inst/n1998 ), .I1(\edb_top_inst/la0/la_trig_pos[14] ), 
            .I2(\edb_top_inst/n2024 ), .I3(\edb_top_inst/la0/la_trig_pos[13] ), 
            .O(\edb_top_inst/n2025 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9ffc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3182 .LUTMASK = 16'h9ffc;
    EFX_LUT4 \edb_top_inst/LUT__3183  (.I0(\edb_top_inst/n1984 ), .I1(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[4] ), .I3(\edb_top_inst/n1981 ), 
            .O(\edb_top_inst/n2026 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3183 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__3184  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n1992 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[8] ), .O(\edb_top_inst/n2027 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf20d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3184 .LUTMASK = 16'hf20d;
    EFX_LUT4 \edb_top_inst/LUT__3185  (.I0(\edb_top_inst/n1989 ), .I1(\edb_top_inst/n1981 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n2028 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b4b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3185 .LUTMASK = 16'h4b4b;
    EFX_LUT4 \edb_top_inst/LUT__3186  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/n2001 ), .I2(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I3(\edb_top_inst/n1982 ), .O(\edb_top_inst/n2029 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb57, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3186 .LUTMASK = 16'heb57;
    EFX_LUT4 \edb_top_inst/LUT__3187  (.I0(\edb_top_inst/n2026 ), .I1(\edb_top_inst/n2028 ), 
            .I2(\edb_top_inst/n2029 ), .I3(\edb_top_inst/n2027 ), .O(\edb_top_inst/n2030 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3187 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3188  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n1986 ), .I2(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n2031 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbff0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3188 .LUTMASK = 16'hbff0;
    EFX_LUT4 \edb_top_inst/LUT__3189  (.I0(\edb_top_inst/n1979 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n2032 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3189 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__3190  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/n1987 ), 
            .I3(\edb_top_inst/n1996 ), .O(\edb_top_inst/n2033 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1428, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3190 .LUTMASK = 16'h1428;
    EFX_LUT4 \edb_top_inst/LUT__3191  (.I0(\edb_top_inst/n2031 ), .I1(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I2(\edb_top_inst/n2032 ), .I3(\edb_top_inst/n2033 ), .O(\edb_top_inst/n2034 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3191 .LUTMASK = 16'h1400;
    EFX_LUT4 \edb_top_inst/LUT__3192  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n2016 ), .I2(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[12] ), .O(\edb_top_inst/n2035 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4fbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3192 .LUTMASK = 16'h4fbb;
    EFX_LUT4 \edb_top_inst/LUT__3193  (.I0(\edb_top_inst/n1981 ), .I1(\edb_top_inst/n1979 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[2] ), .O(\edb_top_inst/n2036 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3193 .LUTMASK = 16'h8787;
    EFX_LUT4 \edb_top_inst/LUT__3194  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .I2(\edb_top_inst/la0/la_trig_pos[16] ), 
            .O(\edb_top_inst/n2037 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3194 .LUTMASK = 16'h8787;
    EFX_LUT4 \edb_top_inst/LUT__3195  (.I0(\edb_top_inst/n1981 ), .I1(\edb_top_inst/n1986 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[1] ), .I3(\edb_top_inst/n2037 ), 
            .O(\edb_top_inst/n2038 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3195 .LUTMASK = 16'h7800;
    EFX_LUT4 \edb_top_inst/LUT__3196  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/n2035 ), .I2(\edb_top_inst/n2036 ), .I3(\edb_top_inst/n2038 ), 
            .O(\edb_top_inst/n2039 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3196 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3197  (.I0(\edb_top_inst/n2025 ), .I1(\edb_top_inst/n2030 ), 
            .I2(\edb_top_inst/n2034 ), .I3(\edb_top_inst/n2039 ), .O(\edb_top_inst/n2040 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3197 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3198  (.I0(\edb_top_inst/n2040 ), .I1(\edb_top_inst/n2003 ), 
            .I2(\edb_top_inst/n2014 ), .I3(\edb_top_inst/n2023 ), .O(\edb_top_inst/n2041 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3198 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3199  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .I2(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n2042 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3199 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3200  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/la0/la_trig_pos[6] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[7] ), .O(\edb_top_inst/n2043 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3200 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3201  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[9] ), .I2(\edb_top_inst/n2042 ), 
            .I3(\edb_top_inst/n2043 ), .O(\edb_top_inst/n2044 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3201 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3202  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[14] ), .I2(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[16] ), .O(\edb_top_inst/n2045 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3202 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3203  (.I0(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[11] ), .I2(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I3(\edb_top_inst/n2045 ), .O(\edb_top_inst/n2046 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3203 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3204  (.I0(\edb_top_inst/n2044 ), .I1(\edb_top_inst/n2046 ), 
            .O(\edb_top_inst/n2047 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3204 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3205  (.I0(\edb_top_inst/la0/la_num_trigger[6] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[7] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .O(\edb_top_inst/n2048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3205 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__3206  (.I0(\edb_top_inst/la0/la_num_trigger[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .O(\edb_top_inst/n2049 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3206 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3207  (.I0(\edb_top_inst/la0/la_num_trigger[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .O(\edb_top_inst/n2050 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3207 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3208  (.I0(\edb_top_inst/n2048 ), .I1(\edb_top_inst/n2049 ), 
            .I2(\edb_top_inst/la0/la_num_trigger[5] ), .I3(\edb_top_inst/n2050 ), 
            .O(\edb_top_inst/n2051 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h333a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3208 .LUTMASK = 16'h333a;
    EFX_LUT4 \edb_top_inst/LUT__3209  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[3] ), .O(\edb_top_inst/n2052 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3209 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3210  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .I2(\edb_top_inst/n2052 ), 
            .I3(\edb_top_inst/n2050 ), .O(\edb_top_inst/n2053 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd6bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3210 .LUTMASK = 16'hd6bf;
    EFX_LUT4 \edb_top_inst/LUT__3211  (.I0(\edb_top_inst/n2050 ), .I1(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I2(\edb_top_inst/n2053 ), .I3(\edb_top_inst/n2051 ), .O(\edb_top_inst/n2054 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3211 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__3212  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[5] ), .I2(\edb_top_inst/la0/la_num_trigger[6] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[7] ), .O(\edb_top_inst/n2055 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3212 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3213  (.I0(\edb_top_inst/la0/la_num_trigger[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), .O(\edb_top_inst/n2056 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3213 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3214  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/n2052 ), .I2(\edb_top_inst/n2055 ), .I3(\edb_top_inst/n2056 ), 
            .O(\edb_top_inst/n2057 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3214 .LUTMASK = 16'hbf40;
    EFX_LUT4 \edb_top_inst/LUT__3215  (.I0(\edb_top_inst/la0/la_num_trigger[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .O(\edb_top_inst/n2058 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3215 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3216  (.I0(\edb_top_inst/la0/la_num_trigger[13] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[14] ), .I2(\edb_top_inst/la0/la_num_trigger[15] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[16] ), .O(\edb_top_inst/n2059 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3216 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3217  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/n2058 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I3(\edb_top_inst/n2059 ), .O(\edb_top_inst/n2060 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3217 .LUTMASK = 16'h1800;
    EFX_LUT4 \edb_top_inst/LUT__3218  (.I0(\edb_top_inst/n2052 ), .I1(\edb_top_inst/n2055 ), 
            .I2(\edb_top_inst/la0/la_num_trigger[8] ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .O(\edb_top_inst/n2061 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7887, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3218 .LUTMASK = 16'h7887;
    EFX_LUT4 \edb_top_inst/LUT__3219  (.I0(\edb_top_inst/la0/la_num_trigger[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .O(\edb_top_inst/n2062 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3219 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3220  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .O(\edb_top_inst/n2063 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3220 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3221  (.I0(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I1(\edb_top_inst/n2062 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I3(\edb_top_inst/n2063 ), .O(\edb_top_inst/n2064 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3221 .LUTMASK = 16'he77b;
    EFX_LUT4 \edb_top_inst/LUT__3222  (.I0(\edb_top_inst/n2064 ), .I1(\edb_top_inst/n2060 ), 
            .I2(\edb_top_inst/n2061 ), .I3(\edb_top_inst/n2057 ), .O(\edb_top_inst/n2065 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3222 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3223  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[9] ), .I2(\edb_top_inst/n2052 ), 
            .I3(\edb_top_inst/n2055 ), .O(\edb_top_inst/n2066 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3223 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3224  (.I0(\edb_top_inst/la0/la_num_trigger[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), .O(\edb_top_inst/n2067 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3224 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3225  (.I0(\edb_top_inst/n2066 ), .I1(\edb_top_inst/la0/la_num_trigger[10] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), .I3(\edb_top_inst/n2067 ), 
            .O(\edb_top_inst/n2068 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb6df, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3225 .LUTMASK = 16'hb6df;
    EFX_LUT4 \edb_top_inst/LUT__3226  (.I0(\edb_top_inst/n2067 ), .I1(\edb_top_inst/la0/la_num_trigger[11] ), 
            .I2(\edb_top_inst/n2066 ), .I3(\edb_top_inst/la0/la_num_trigger[12] ), 
            .O(\edb_top_inst/n2069 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef15, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3226 .LUTMASK = 16'hef15;
    EFX_LUT4 \edb_top_inst/LUT__3227  (.I0(\edb_top_inst/n2068 ), .I1(\edb_top_inst/n2069 ), 
            .I2(\edb_top_inst/n2054 ), .I3(\edb_top_inst/n2065 ), .O(\edb_top_inst/n2070 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3227 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3228  (.I0(\edb_top_inst/n2047 ), .I1(\edb_top_inst/n2070 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2071 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3228 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3229  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n1984 ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[12] ), .O(\edb_top_inst/n2072 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf807, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3229 .LUTMASK = 16'hf807;
    EFX_LUT4 \edb_top_inst/LUT__3230  (.I0(\edb_top_inst/n1995 ), .I1(\edb_top_inst/n1996 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[0] ), .O(\edb_top_inst/n2073 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8787, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3230 .LUTMASK = 16'h8787;
    EFX_LUT4 \edb_top_inst/LUT__3231  (.I0(\edb_top_inst/n2073 ), .I1(\edb_top_inst/n2036 ), 
            .I2(\edb_top_inst/n2072 ), .I3(\edb_top_inst/n2038 ), .O(\edb_top_inst/n2074 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3231 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3232  (.I0(\edb_top_inst/n2025 ), .I1(\edb_top_inst/n2030 ), 
            .I2(\edb_top_inst/n2034 ), .I3(\edb_top_inst/n2074 ), .O(\edb_top_inst/n2075 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3232 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3233  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n2076 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3233 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3234  (.I0(\edb_top_inst/n2075 ), .I1(\edb_top_inst/la0/la_stop_trig ), 
            .I2(\edb_top_inst/n1978 ), .I3(\edb_top_inst/n2076 ), .O(\edb_top_inst/n2077 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3234 .LUTMASK = 16'h3a00;
    EFX_LUT4 \edb_top_inst/LUT__3235  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[10] ), .I2(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[12] ), .O(\edb_top_inst/n2078 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf5dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3235 .LUTMASK = 16'hf5dc;
    EFX_LUT4 \edb_top_inst/LUT__3236  (.I0(\edb_top_inst/n2044 ), .I1(\edb_top_inst/n2078 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[12] ), .I3(\edb_top_inst/n2045 ), 
            .O(\edb_top_inst/n2079 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3236 .LUTMASK = 16'h3d00;
    EFX_LUT4 \edb_top_inst/LUT__3237  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I2(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n2080 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3237 .LUTMASK = 16'hbed7;
    EFX_LUT4 \edb_top_inst/LUT__3238  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[6] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[7] ), .O(\edb_top_inst/n2081 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3238 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3239  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n2082 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3239 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3240  (.I0(\edb_top_inst/n2080 ), .I1(\edb_top_inst/n2081 ), 
            .I2(\edb_top_inst/n2042 ), .I3(\edb_top_inst/n2082 ), .O(\edb_top_inst/n2083 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha333, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3240 .LUTMASK = 16'ha333;
    EFX_LUT4 \edb_top_inst/LUT__3241  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[9] ), .O(\edb_top_inst/n2084 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb00b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3241 .LUTMASK = 16'hb00b;
    EFX_LUT4 \edb_top_inst/LUT__3242  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), .O(\edb_top_inst/n2085 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3242 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3243  (.I0(\edb_top_inst/n2084 ), .I1(\edb_top_inst/n2085 ), 
            .I2(\edb_top_inst/n2042 ), .I3(\edb_top_inst/n2043 ), .O(\edb_top_inst/n2086 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5333, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3243 .LUTMASK = 16'h5333;
    EFX_LUT4 \edb_top_inst/LUT__3244  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I2(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .O(\edb_top_inst/n2087 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3244 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__3245  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .O(\edb_top_inst/n2088 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3245 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3246  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n2089 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3246 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3247  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[2] ), .I2(\edb_top_inst/n2088 ), 
            .I3(\edb_top_inst/n2089 ), .O(\edb_top_inst/n2090 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb6df, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3247 .LUTMASK = 16'hb6df;
    EFX_LUT4 \edb_top_inst/LUT__3248  (.I0(\edb_top_inst/n2083 ), .I1(\edb_top_inst/n2087 ), 
            .I2(\edb_top_inst/n2090 ), .I3(\edb_top_inst/n2086 ), .O(\edb_top_inst/n2091 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3248 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3249  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), .I2(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[4] ), .O(\edb_top_inst/n2092 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbed7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3249 .LUTMASK = 16'hbed7;
    EFX_LUT4 \edb_top_inst/LUT__3250  (.I0(\edb_top_inst/n2085 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[9] ), .O(\edb_top_inst/n2093 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3250 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__3251  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[4] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n2094 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3251 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3252  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .O(\edb_top_inst/n2095 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3252 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3253  (.I0(\edb_top_inst/n2043 ), .I1(\edb_top_inst/n2094 ), 
            .I2(\edb_top_inst/n2042 ), .I3(\edb_top_inst/n2095 ), .O(\edb_top_inst/n2096 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5f03, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3253 .LUTMASK = 16'h5f03;
    EFX_LUT4 \edb_top_inst/LUT__3254  (.I0(\edb_top_inst/n2092 ), .I1(\edb_top_inst/n2042 ), 
            .I2(\edb_top_inst/n2093 ), .I3(\edb_top_inst/n2096 ), .O(\edb_top_inst/n2097 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3254 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3255  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[11] ), .O(\edb_top_inst/n2098 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3255 .LUTMASK = 16'h9999;
    EFX_LUT4 \edb_top_inst/LUT__3256  (.I0(\edb_top_inst/n2098 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I2(\edb_top_inst/n2044 ), .I3(\edb_top_inst/la0/la_trig_pos[10] ), 
            .O(\edb_top_inst/n2099 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd73d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3256 .LUTMASK = 16'hd73d;
    EFX_LUT4 \edb_top_inst/LUT__3257  (.I0(\edb_top_inst/n2099 ), .I1(\edb_top_inst/n2091 ), 
            .I2(\edb_top_inst/n2097 ), .I3(\edb_top_inst/n2079 ), .O(\edb_top_inst/n2100 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3257 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3258  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n2101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3258 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3259  (.I0(\edb_top_inst/n2101 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n2047 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2102 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00fe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3259 .LUTMASK = 16'h00fe;
    EFX_LUT4 \edb_top_inst/LUT__3260  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n2103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3260 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3261  (.I0(\edb_top_inst/n2100 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n2102 ), .I3(\edb_top_inst/n2103 ), .O(\edb_top_inst/n2104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3261 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__3262  (.I0(\edb_top_inst/n2071 ), .I1(\edb_top_inst/n2041 ), 
            .I2(\edb_top_inst/n2077 ), .I3(\edb_top_inst/n2104 ), .O(\edb_top_inst/n2105 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3262 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__3263  (.I0(\edb_top_inst/n2100 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I2(\edb_top_inst/n2005 ), .O(\edb_top_inst/n2106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3263 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3264  (.I0(\edb_top_inst/n2006 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n2105 ), .I3(\edb_top_inst/n2106 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3264 .LUTMASK = 16'hfff4;
    EFX_LUT4 \edb_top_inst/LUT__3265  (.I0(\edb_top_inst/n1801 ), .I1(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/la0/la_biu_inst/n350 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3265 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3266  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/n1251 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3266 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3267  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), .I2(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q ), 
            .I3(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3267 .LUTMASK = 16'h00be;
    EFX_LUT4 \edb_top_inst/LUT__3268  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .I2(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .O(\edb_top_inst/ceg_net351 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3268 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3269  (.I0(\edb_top_inst/n1978 ), .I1(\edb_top_inst/n2075 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/n2005 ), 
            .O(\edb_top_inst/n2107 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3269 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__3270  (.I0(\edb_top_inst/n1978 ), .I1(\edb_top_inst/n2070 ), 
            .I2(\edb_top_inst/n2003 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3270 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__3271  (.I0(\edb_top_inst/n2047 ), .I1(\edb_top_inst/n2070 ), 
            .O(\edb_top_inst/n2109 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3271 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3272  (.I0(\edb_top_inst/n2041 ), .I1(\edb_top_inst/n2109 ), 
            .I2(\edb_top_inst/n2108 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n2110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3272 .LUTMASK = 16'h0fbb;
    EFX_LUT4 \edb_top_inst/LUT__3273  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n2110 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I3(\edb_top_inst/n2107 ), .O(\edb_top_inst/la0/la_biu_inst/n1236 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3273 .LUTMASK = 16'h8700;
    EFX_LUT4 \edb_top_inst/LUT__3274  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/n7224 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3274 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3275  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/n2103 ), .O(\edb_top_inst/n2111 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3275 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3276  (.I0(\edb_top_inst/n1872 ), .I1(\edb_top_inst/n2109 ), 
            .I2(\edb_top_inst/n2111 ), .O(\edb_top_inst/n2112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3276 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3277  (.I0(\edb_top_inst/n2070 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n2113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3277 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3278  (.I0(\edb_top_inst/n1978 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n2114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3278 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3279  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n2115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3279 .LUTMASK = 16'hfa3f;
    EFX_LUT4 \edb_top_inst/LUT__3280  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/n2003 ), .I2(\edb_top_inst/n2114 ), .I3(\edb_top_inst/n2115 ), 
            .O(\edb_top_inst/n2116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3280 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__3281  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n2113 ), .I2(\edb_top_inst/n2116 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n2117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3281 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3282  (.I0(\edb_top_inst/n2075 ), .I1(\edb_top_inst/n2070 ), 
            .I2(\edb_top_inst/la0/la_stop_trig ), .I3(\edb_top_inst/n1978 ), 
            .O(\edb_top_inst/n2118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3282 .LUTMASK = 16'h0fbb;
    EFX_LUT4 \edb_top_inst/LUT__3283  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3283 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3284  (.I0(\edb_top_inst/n2118 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I2(\edb_top_inst/n2119 ), .O(\edb_top_inst/n2120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3284 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__3285  (.I0(\edb_top_inst/n2112 ), .I1(\edb_top_inst/n2041 ), 
            .I2(\edb_top_inst/n2117 ), .I3(\edb_top_inst/n2120 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3285 .LUTMASK = 16'hfff2;
    EFX_LUT4 \edb_top_inst/LUT__3286  (.I0(\edb_top_inst/la0/la_stop_trig ), 
            .I1(\edb_top_inst/n2075 ), .I2(\edb_top_inst/n2070 ), .I3(\edb_top_inst/n1978 ), 
            .O(\edb_top_inst/n2121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h55c3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3286 .LUTMASK = 16'h55c3;
    EFX_LUT4 \edb_top_inst/LUT__3287  (.I0(\edb_top_inst/n2070 ), .I1(\edb_top_inst/n2047 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n2122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3287 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__3288  (.I0(\edb_top_inst/n2041 ), .I1(\edb_top_inst/n2122 ), 
            .I2(\edb_top_inst/n2121 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n2123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3288 .LUTMASK = 16'hbbb0;
    EFX_LUT4 \edb_top_inst/LUT__3289  (.I0(\edb_top_inst/n2101 ), .I1(\edb_top_inst/n2047 ), 
            .I2(\edb_top_inst/n1872 ), .I3(\edb_top_inst/n2005 ), .O(\edb_top_inst/n2124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3289 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3290  (.I0(\edb_top_inst/n2005 ), .I1(\edb_top_inst/n2116 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/n2100 ), 
            .O(\edb_top_inst/n2125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h133f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3290 .LUTMASK = 16'h133f;
    EFX_LUT4 \edb_top_inst/LUT__3291  (.I0(\edb_top_inst/n2111 ), .I1(\edb_top_inst/n2123 ), 
            .I2(\edb_top_inst/n2124 ), .I3(\edb_top_inst/n2125 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3291 .LUTMASK = 16'hf8ff;
    EFX_LUT4 \edb_top_inst/LUT__3292  (.I0(\edb_top_inst/la0/la_biu_inst/n350 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ), .I2(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
            .O(\edb_top_inst/ceg_net348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3292 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__3293  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3293 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3294  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n2119 ), .I2(\edb_top_inst/n1978 ), .O(\edb_top_inst/la0/la_biu_inst/n1993 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfbf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3294 .LUTMASK = 16'hbfbf;
    EFX_LUT4 \edb_top_inst/LUT__3295  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/la0/la_biu_inst/fifo_push )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05fc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3295 .LUTMASK = 16'h05fc;
    EFX_LUT4 \edb_top_inst/LUT__3296  (.I0(\edb_top_inst/la0/la_biu_inst/n1993 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_push ), .O(\edb_top_inst/n2126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3296 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3297  (.I0(\edb_top_inst/n2126 ), .I1(\edb_top_inst/n2003 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3297 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3298  (.I0(\edb_top_inst/n2005 ), .I1(\edb_top_inst/n1872 ), 
            .I2(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_rstn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3298 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3299  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3299 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3300  (.I0(\edb_top_inst/n2126 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
            .O(\edb_top_inst/ceg_net355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3300 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3301  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ), 
            .I1(\edb_top_inst/n1873 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3301 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3302  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[15] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3302 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3303  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[16] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3303 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3304  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[17] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3304 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3305  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[18] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3305 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3306  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[19] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3306 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3307  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[20] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3307 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3308  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[21] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3308 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3309  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[22] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3309 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3310  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[23] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3310 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3311  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[24] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3311 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3312  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[25] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3312 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3313  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[26] ), .I2(\edb_top_inst/n1873 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3313 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3314  (.I0(\edb_top_inst/n1995 ), .I1(\edb_top_inst/n1996 ), 
            .O(\edb_top_inst/n2127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3314 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3315  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .I1(\edb_top_inst/n2017 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I3(\edb_top_inst/n2127 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3315 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__3316  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/n2011 ), .O(\edb_top_inst/n2128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3316 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3317  (.I0(\edb_top_inst/n1984 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n2129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3317 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3318  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .I3(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3318 .LUTMASK = 16'h0c0a;
    EFX_LUT4 \edb_top_inst/LUT__3319  (.I0(\edb_top_inst/n1996 ), .I1(\edb_top_inst/n2130 ), 
            .O(\edb_top_inst/n2131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3319 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3320  (.I0(\edb_top_inst/n2128 ), .I1(\edb_top_inst/n2129 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I3(\edb_top_inst/n2131 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3320 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3321  (.I0(\edb_top_inst/n1984 ), .I1(\edb_top_inst/n1999 ), 
            .O(\edb_top_inst/n2132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3321 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3322  (.I0(\edb_top_inst/n1979 ), .I1(\edb_top_inst/n1981 ), 
            .I2(\edb_top_inst/n2132 ), .O(\edb_top_inst/n2133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3322 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__3323  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3323 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3324  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/n2134 ), 
            .I3(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3324 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3325  (.I0(\edb_top_inst/n2135 ), .I1(\edb_top_inst/n1996 ), 
            .I2(\edb_top_inst/n2133 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3325 .LUTMASK = 16'h4f44;
    EFX_LUT4 \edb_top_inst/LUT__3326  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3326 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3327  (.I0(\edb_top_inst/n2136 ), .I1(\edb_top_inst/n2134 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3327 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3328  (.I0(\edb_top_inst/n2137 ), .I1(\edb_top_inst/n1996 ), 
            .O(\edb_top_inst/n2138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3328 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3329  (.I0(\edb_top_inst/n2011 ), .I1(\edb_top_inst/n2129 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I3(\edb_top_inst/n2138 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3329 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3330  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n2015 ), .O(\edb_top_inst/n2139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3330 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3331  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I1(\edb_top_inst/n1995 ), .O(\edb_top_inst/n2140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3331 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3332  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3332 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3333  (.I0(\edb_top_inst/n2141 ), .I1(\edb_top_inst/n2136 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3333 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3334  (.I0(\edb_top_inst/n2142 ), .I1(\edb_top_inst/n2140 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n1981 ), 
            .O(\edb_top_inst/n2143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3334 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__3335  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I1(\edb_top_inst/n2139 ), .I2(\edb_top_inst/n2143 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3335 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3336  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .I3(\edb_top_inst/n2139 ), .O(\edb_top_inst/n2144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3336 .LUTMASK = 16'hbf00;
    EFX_LUT4 \edb_top_inst/LUT__3337  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3337 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3338  (.I0(\edb_top_inst/n2145 ), .I1(\edb_top_inst/n2141 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3338 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3339  (.I0(\edb_top_inst/n2146 ), .I1(\edb_top_inst/n2130 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n1981 ), 
            .O(\edb_top_inst/n2147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3339 .LUTMASK = 16'hc500;
    EFX_LUT4 \edb_top_inst/LUT__3340  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I1(\edb_top_inst/n2144 ), .I2(\edb_top_inst/n2147 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3340 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3341  (.I0(\edb_top_inst/n1998 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n2144 ), .O(\edb_top_inst/n2148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3341 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3342  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3342 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3343  (.I0(\edb_top_inst/n2149 ), .I1(\edb_top_inst/n2145 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3343 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3344  (.I0(\edb_top_inst/n2150 ), .I1(\edb_top_inst/n2135 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n1981 ), 
            .O(\edb_top_inst/n2151 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3344 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__3345  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I1(\edb_top_inst/n2148 ), .I2(\edb_top_inst/n2151 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3345 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3346  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3346 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3347  (.I0(\edb_top_inst/n2152 ), .I1(\edb_top_inst/n2149 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2153 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3347 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3348  (.I0(\edb_top_inst/n2153 ), .I1(\edb_top_inst/n2137 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n1981 ), 
            .O(\edb_top_inst/n2154 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3348 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__3349  (.I0(\edb_top_inst/n2132 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I2(\edb_top_inst/n2154 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3349 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3350  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2155 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3350 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3351  (.I0(\edb_top_inst/n2155 ), .I1(\edb_top_inst/n2152 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3351 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3352  (.I0(\edb_top_inst/n2156 ), .I1(\edb_top_inst/n2140 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n2157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf30a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3352 .LUTMASK = 16'hf30a;
    EFX_LUT4 \edb_top_inst/LUT__3353  (.I0(\edb_top_inst/n2142 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n2157 ), 
            .O(\edb_top_inst/n2158 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3353 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3354  (.I0(\edb_top_inst/n1992 ), .I1(\edb_top_inst/n2132 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I3(\edb_top_inst/n2158 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3354 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3355  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n2159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3355 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__3356  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3356 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3357  (.I0(\edb_top_inst/n2160 ), .I1(\edb_top_inst/n2155 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3357 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3358  (.I0(\edb_top_inst/n2161 ), .I1(\edb_top_inst/n2130 ), 
            .I2(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n2162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3358 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__3359  (.I0(\edb_top_inst/n2162 ), .I1(\edb_top_inst/n2146 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n1982 ), 
            .O(\edb_top_inst/n2163 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3359 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__3360  (.I0(\edb_top_inst/n2159 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I2(\edb_top_inst/n2139 ), .I3(\edb_top_inst/n2163 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3360 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3361  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2164 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3361 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3362  (.I0(\edb_top_inst/n2164 ), .I1(\edb_top_inst/n2160 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2165 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3362 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3363  (.I0(\edb_top_inst/n2165 ), .I1(\edb_top_inst/n2150 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n1981 ), 
            .O(\edb_top_inst/n2166 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3363 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__3364  (.I0(\edb_top_inst/n2135 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n1999 ), .I3(\edb_top_inst/n2166 ), .O(\edb_top_inst/n2167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3364 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__3365  (.I0(\edb_top_inst/n1979 ), .I1(\edb_top_inst/n2132 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] ), 
            .I3(\edb_top_inst/n2167 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3365 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__3366  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n1995 ), .O(\edb_top_inst/n2168 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3366 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3367  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3367 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__3368  (.I0(\edb_top_inst/n2169 ), .I1(\edb_top_inst/n2164 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2170 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3368 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3369  (.I0(\edb_top_inst/n2170 ), .I1(\edb_top_inst/n2153 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n1981 ), 
            .O(\edb_top_inst/n2171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3369 .LUTMASK = 16'h3500;
    EFX_LUT4 \edb_top_inst/LUT__3370  (.I0(\edb_top_inst/n2137 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n1999 ), .I3(\edb_top_inst/n2171 ), .O(\edb_top_inst/n2172 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3370 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__3371  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] ), 
            .I1(\edb_top_inst/n1999 ), .I2(\edb_top_inst/n2168 ), .I3(\edb_top_inst/n2172 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h80ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3371 .LUTMASK = 16'h80ff;
    EFX_LUT4 \edb_top_inst/LUT__3372  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .I1(\edb_top_inst/n2017 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I3(\edb_top_inst/n2127 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3372 .LUTMASK = 16'hf888;
    EFX_LUT4 \edb_top_inst/LUT__3373  (.I0(\edb_top_inst/n2128 ), .I1(\edb_top_inst/n2129 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I3(\edb_top_inst/n2131 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3373 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3374  (.I0(\edb_top_inst/n2135 ), .I1(\edb_top_inst/n1996 ), 
            .I2(\edb_top_inst/n2133 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3374 .LUTMASK = 16'h4f44;
    EFX_LUT4 \edb_top_inst/LUT__3375  (.I0(\edb_top_inst/n2011 ), .I1(\edb_top_inst/n2129 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I3(\edb_top_inst/n2138 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3375 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3376  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I1(\edb_top_inst/n2139 ), .I2(\edb_top_inst/n2143 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3376 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3377  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I1(\edb_top_inst/n2144 ), .I2(\edb_top_inst/n2147 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3377 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3378  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I1(\edb_top_inst/n2148 ), .I2(\edb_top_inst/n2151 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3378 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3379  (.I0(\edb_top_inst/n2132 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I2(\edb_top_inst/n2154 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3379 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3380  (.I0(\edb_top_inst/n1992 ), .I1(\edb_top_inst/n2132 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I3(\edb_top_inst/n2158 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3380 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3381  (.I0(\edb_top_inst/n2159 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I2(\edb_top_inst/n2139 ), .I3(\edb_top_inst/n2163 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3381 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__3382  (.I0(\edb_top_inst/n1979 ), .I1(\edb_top_inst/n2132 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] ), 
            .I3(\edb_top_inst/n2167 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3382 .LUTMASK = 16'h40ff;
    EFX_LUT4 \edb_top_inst/LUT__3383  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] ), 
            .I1(\edb_top_inst/n1999 ), .I2(\edb_top_inst/n2168 ), .I3(\edb_top_inst/n2172 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h80ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3383 .LUTMASK = 16'h80ff;
    EFX_LUT4 \edb_top_inst/LUT__3384  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .I2(\edb_top_inst/la0/module_state[0] ), 
            .I3(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n2173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcc53, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3384 .LUTMASK = 16'hcc53;
    EFX_LUT4 \edb_top_inst/LUT__3385  (.I0(\edb_top_inst/n2173 ), .I1(jtag_inst1_UPDATE), 
            .I2(\edb_top_inst/edb_user_dr[81] ), .I3(jtag_inst1_SEL), .O(\edb_top_inst/debug_hub_inst/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3385 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3386  (.I0(jtag_inst1_SEL), .I1(jtag_inst1_SHIFT), 
            .O(\edb_top_inst/debug_hub_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3386 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3387  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[1] ), .O(\edb_top_inst/n1711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3387 .LUTMASK = 16'h1000;
    EFX_ADD \edb_top_inst/la0/add_91/i1  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/n969 ), .CI(1'b0), .O(\edb_top_inst/n34 ), 
            .CO(\edb_top_inst/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i2  (.I0(\edb_top_inst/la0/bit_count[1] ), 
            .I1(\edb_top_inst/la0/bit_count[0] ), .CI(1'b0), .O(\edb_top_inst/n36 ), 
            .CO(\edb_top_inst/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/add_100/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .CI(1'b0), 
            .O(\edb_top_inst/n297 ), .CO(\edb_top_inst/n298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/n426 ), .CO(\edb_top_inst/n427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/n428 ), .CO(\edb_top_inst/n429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .CI(1'b0), 
            .O(\edb_top_inst/n432 ), .CO(\edb_top_inst/n433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[0] ), .CI(1'b0), .O(\edb_top_inst/n434 ), 
            .CO(\edb_top_inst/n435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13  (.I0(\edb_top_inst/la0/la_sample_cnt[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n613 ), .O(\edb_top_inst/n590 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12  (.I0(\edb_top_inst/la0/la_sample_cnt[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n615 ), .O(\edb_top_inst/n612 ), 
            .CO(\edb_top_inst/n613 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n617 ), .O(\edb_top_inst/n614 ), 
            .CO(\edb_top_inst/n615 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n619 ), .O(\edb_top_inst/n616 ), 
            .CO(\edb_top_inst/n617 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n621 ), .O(\edb_top_inst/n618 ), 
            .CO(\edb_top_inst/n619 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n623 ), .O(\edb_top_inst/n620 ), 
            .CO(\edb_top_inst/n621 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n625 ), .O(\edb_top_inst/n622 ), 
            .CO(\edb_top_inst/n623 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n627 ), .O(\edb_top_inst/n624 ), 
            .CO(\edb_top_inst/n625 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n629 ), .O(\edb_top_inst/n626 ), 
            .CO(\edb_top_inst/n627 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n631 ), .O(\edb_top_inst/n628 ), 
            .CO(\edb_top_inst/n629 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n435 ), .O(\edb_top_inst/n630 ), 
            .CO(\edb_top_inst/n631 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4635)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n634 ), .O(\edb_top_inst/n632 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n636 ), .O(\edb_top_inst/n633 ), 
            .CO(\edb_top_inst/n634 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n638 ), .O(\edb_top_inst/n635 ), 
            .CO(\edb_top_inst/n636 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n640 ), .O(\edb_top_inst/n637 ), 
            .CO(\edb_top_inst/n638 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n642 ), .O(\edb_top_inst/n639 ), 
            .CO(\edb_top_inst/n640 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n644 ), .O(\edb_top_inst/n641 ), 
            .CO(\edb_top_inst/n642 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n646 ), .O(\edb_top_inst/n643 ), 
            .CO(\edb_top_inst/n644 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n648 ), .O(\edb_top_inst/n645 ), 
            .CO(\edb_top_inst/n646 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n650 ), .O(\edb_top_inst/n647 ), 
            .CO(\edb_top_inst/n648 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n652 ), .O(\edb_top_inst/n649 ), 
            .CO(\edb_top_inst/n650 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n433 ), .O(\edb_top_inst/n651 ), 
            .CO(\edb_top_inst/n652 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4621)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n680 ), .O(\edb_top_inst/n677 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n682 ), .O(\edb_top_inst/n679 ), 
            .CO(\edb_top_inst/n680 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n684 ), .O(\edb_top_inst/n681 ), 
            .CO(\edb_top_inst/n682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n686 ), .O(\edb_top_inst/n683 ), 
            .CO(\edb_top_inst/n684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n688 ), .O(\edb_top_inst/n685 ), 
            .CO(\edb_top_inst/n686 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n690 ), .O(\edb_top_inst/n687 ), 
            .CO(\edb_top_inst/n688 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n692 ), .O(\edb_top_inst/n689 ), 
            .CO(\edb_top_inst/n690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n694 ), .O(\edb_top_inst/n691 ), 
            .CO(\edb_top_inst/n692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n696 ), .O(\edb_top_inst/n693 ), 
            .CO(\edb_top_inst/n694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n429 ), .O(\edb_top_inst/n695 ), 
            .CO(\edb_top_inst/n696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4614)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n731 ), .O(\edb_top_inst/n727 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n733 ), .O(\edb_top_inst/n730 ), 
            .CO(\edb_top_inst/n731 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n735 ), .O(\edb_top_inst/n732 ), 
            .CO(\edb_top_inst/n733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n737 ), .O(\edb_top_inst/n734 ), 
            .CO(\edb_top_inst/n735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n739 ), .O(\edb_top_inst/n736 ), 
            .CO(\edb_top_inst/n737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n741 ), .O(\edb_top_inst/n738 ), 
            .CO(\edb_top_inst/n739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n743 ), .O(\edb_top_inst/n740 ), 
            .CO(\edb_top_inst/n741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n745 ), .O(\edb_top_inst/n742 ), 
            .CO(\edb_top_inst/n743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n747 ), .O(\edb_top_inst/n744 ), 
            .CO(\edb_top_inst/n745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n427 ), .O(\edb_top_inst/n746 ), 
            .CO(\edb_top_inst/n747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4610)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n750 ), .O(\edb_top_inst/n748 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n752 ), .O(\edb_top_inst/n749 ), 
            .CO(\edb_top_inst/n750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n754 ), .O(\edb_top_inst/n751 ), 
            .CO(\edb_top_inst/n752 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n756 ), .O(\edb_top_inst/n753 ), 
            .CO(\edb_top_inst/n754 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n758 ), .O(\edb_top_inst/n755 ), 
            .CO(\edb_top_inst/n756 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n760 ), .O(\edb_top_inst/n757 ), 
            .CO(\edb_top_inst/n758 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n762 ), .O(\edb_top_inst/n759 ), 
            .CO(\edb_top_inst/n760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n764 ), .O(\edb_top_inst/n761 ), 
            .CO(\edb_top_inst/n762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n766 ), .O(\edb_top_inst/n763 ), 
            .CO(\edb_top_inst/n764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n298 ), .O(\edb_top_inst/n765 ), 
            .CO(\edb_top_inst/n766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(4603)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i6  (.I0(\edb_top_inst/la0/bit_count[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n769 ), .O(\edb_top_inst/n767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/add_100/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i5  (.I0(\edb_top_inst/la0/bit_count[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n771 ), .O(\edb_top_inst/n768 ), 
            .CO(\edb_top_inst/n769 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/add_100/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i4  (.I0(\edb_top_inst/la0/bit_count[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n773 ), .O(\edb_top_inst/n770 ), 
            .CO(\edb_top_inst/n771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/add_100/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i3  (.I0(\edb_top_inst/la0/bit_count[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n37 ), .O(\edb_top_inst/n772 ), 
            .CO(\edb_top_inst/n773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3681)
    defparam \edb_top_inst/la0/add_100/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i27  (.I0(\edb_top_inst/la0/address_counter[26] ), 
            .I1(1'b0), .CI(\edb_top_inst/n786 ), .O(\edb_top_inst/n783 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i27 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i26  (.I0(\edb_top_inst/la0/address_counter[25] ), 
            .I1(1'b0), .CI(\edb_top_inst/n788 ), .O(\edb_top_inst/n785 ), 
            .CO(\edb_top_inst/n786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i26 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i25  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/n790 ), .O(\edb_top_inst/n787 ), 
            .CO(\edb_top_inst/n788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i24  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/n792 ), .O(\edb_top_inst/n789 ), 
            .CO(\edb_top_inst/n790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i23  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/n794 ), .O(\edb_top_inst/n791 ), 
            .CO(\edb_top_inst/n792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i22  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/n796 ), .O(\edb_top_inst/n793 ), 
            .CO(\edb_top_inst/n794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i21  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/n798 ), .O(\edb_top_inst/n795 ), 
            .CO(\edb_top_inst/n796 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i20  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/n800 ), .O(\edb_top_inst/n797 ), 
            .CO(\edb_top_inst/n798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i19  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/n802 ), .O(\edb_top_inst/n799 ), 
            .CO(\edb_top_inst/n800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i18  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/n804 ), .O(\edb_top_inst/n801 ), 
            .CO(\edb_top_inst/n802 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i17  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(1'b0), .CI(\edb_top_inst/n806 ), .O(\edb_top_inst/n803 ), 
            .CO(\edb_top_inst/n804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i16  (.I0(\edb_top_inst/la0/address_counter[15] ), 
            .I1(1'b0), .CI(\edb_top_inst/n808 ), .O(\edb_top_inst/n805 ), 
            .CO(\edb_top_inst/n806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i15  (.I0(\edb_top_inst/la0/address_counter[14] ), 
            .I1(1'b0), .CI(\edb_top_inst/n810 ), .O(\edb_top_inst/n807 ), 
            .CO(\edb_top_inst/n808 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i14  (.I0(\edb_top_inst/la0/address_counter[13] ), 
            .I1(1'b0), .CI(\edb_top_inst/n812 ), .O(\edb_top_inst/n809 ), 
            .CO(\edb_top_inst/n810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i13  (.I0(\edb_top_inst/la0/address_counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n814 ), .O(\edb_top_inst/n811 ), 
            .CO(\edb_top_inst/n812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i12  (.I0(\edb_top_inst/la0/address_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n816 ), .O(\edb_top_inst/n813 ), 
            .CO(\edb_top_inst/n814 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i11  (.I0(\edb_top_inst/la0/address_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n818 ), .O(\edb_top_inst/n815 ), 
            .CO(\edb_top_inst/n816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i10  (.I0(\edb_top_inst/la0/address_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n820 ), .O(\edb_top_inst/n817 ), 
            .CO(\edb_top_inst/n818 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i9  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n822 ), .O(\edb_top_inst/n819 ), 
            .CO(\edb_top_inst/n820 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i8  (.I0(\edb_top_inst/la0/address_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n824 ), .O(\edb_top_inst/n821 ), 
            .CO(\edb_top_inst/n822 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i7  (.I0(\edb_top_inst/la0/address_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n826 ), .O(\edb_top_inst/n823 ), 
            .CO(\edb_top_inst/n824 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i6  (.I0(\edb_top_inst/la0/address_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n828 ), .O(\edb_top_inst/n825 ), 
            .CO(\edb_top_inst/n826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i5  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n830 ), .O(\edb_top_inst/n827 ), 
            .CO(\edb_top_inst/n828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i4  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/n1705 ), .CI(\edb_top_inst/n832 ), .O(\edb_top_inst/n829 ), 
            .CO(\edb_top_inst/n830 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i3  (.I0(\edb_top_inst/la0/address_counter[2] ), 
            .I1(\edb_top_inst/n1708 ), .CI(\edb_top_inst/n834 ), .O(\edb_top_inst/n831 ), 
            .CO(\edb_top_inst/n832 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i2  (.I0(\edb_top_inst/la0/address_counter[1] ), 
            .I1(\edb_top_inst/n1711 ), .CI(\edb_top_inst/n35 ), .O(\edb_top_inst/n833 ), 
            .CO(\edb_top_inst/n834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3654)
    defparam \edb_top_inst/la0/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i12  (.I0(\edb_top_inst/la0/address_counter[26] ), 
            .I1(1'b0), .CI(\edb_top_inst/n847 ), .O(\edb_top_inst/n844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i11  (.I0(\edb_top_inst/la0/address_counter[25] ), 
            .I1(1'b0), .CI(\edb_top_inst/n849 ), .O(\edb_top_inst/n846 ), 
            .CO(\edb_top_inst/n847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i10  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/n851 ), .O(\edb_top_inst/n848 ), 
            .CO(\edb_top_inst/n849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i9  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/n853 ), .O(\edb_top_inst/n850 ), 
            .CO(\edb_top_inst/n851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i8  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/n855 ), .O(\edb_top_inst/n852 ), 
            .CO(\edb_top_inst/n853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i7  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/n857 ), .O(\edb_top_inst/n854 ), 
            .CO(\edb_top_inst/n855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i6  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/n862 ), .O(\edb_top_inst/n856 ), 
            .CO(\edb_top_inst/n857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i5  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/n864 ), .O(\edb_top_inst/n861 ), 
            .CO(\edb_top_inst/n862 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i4  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/n866 ), .O(\edb_top_inst/n863 ), 
            .CO(\edb_top_inst/n864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i3  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/n868 ), .O(\edb_top_inst/n865 ), 
            .CO(\edb_top_inst/n866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i2  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(\edb_top_inst/la0/address_counter[15] ), .CI(1'b0), .O(\edb_top_inst/n867 ), 
            .CO(\edb_top_inst/n868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(3653)
    defparam \edb_top_inst/la0/add_90/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i2 .I1_POLARITY = 1'b1;
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2090), .WDATA({\cmos_frame_Gray[0] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n105 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2104), .WDATA({\cmos_frame_Gray[2] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n98 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2090), .WDATA({\cmos_frame_Gray[2] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n99 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2090), .WDATA({\cmos_frame_Gray[1] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n102 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2104), .WDATA({\cmos_frame_Gray[0] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n104 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2090), .WDATA({\cmos_frame_Gray[3] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n96 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2090), .WDATA({\cmos_frame_Gray[4] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n93 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2090), .WDATA({\cmos_frame_Gray[5] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n90 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2090), .WDATA({\cmos_frame_Gray[6] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n87 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2090), .WDATA({\cmos_frame_Gray[7] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n84 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2104), .WDATA({\cmos_frame_Gray[1] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n101 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2104), .WDATA({\cmos_frame_Gray[3] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n95 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2104), .WDATA({\cmos_frame_Gray[4] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n92 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2104), .WDATA({\cmos_frame_Gray[5] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n89 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2104), .WDATA({\cmos_frame_Gray[6] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n86 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2104), .WDATA({\cmos_frame_Gray[7] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n83 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[6] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_1=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_2=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_3=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_4=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_5=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_6=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_7=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_0 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_1 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_2 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_3 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_4 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_5 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_6 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_7 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[1] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_1=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_2=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_3=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_4=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_5=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_6=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_7=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_0 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_1 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_2 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_3 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_4 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_5 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_6 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_7 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[1] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_1=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_2=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_3=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_4=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_5=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_6=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_7=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_0 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_1 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_2 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_3 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_4 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_5 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_6 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_7 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[1] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_1=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_2=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_3=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_4=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_5=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_6=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_7=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_0 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_1 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_2 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_3 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_4 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_5 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_6 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_7 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[1] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_1=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_2=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_3=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_4=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_5=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_6=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_7=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_0 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_1 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_2 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_3 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_4 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_5 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_6 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_7 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[5] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_1=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_2=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_3=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_4=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_5=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_6=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_7=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_0 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_1 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_2 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_3 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_4 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_5 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_6 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_7 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[7] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_1=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_2=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_3=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_4=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_5=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_6=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_7=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_0 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_1 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_2 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_3 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_4 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_5 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_6 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_7 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[4] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_1=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_2=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_3=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_4=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_5=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_6=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_7=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_0 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_1 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_2 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_3 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_4 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_5 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_6 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_7 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[2] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_1=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_2=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_3=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_4=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_5=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_6=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_7=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_0 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_1 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_2 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_3 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_4 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_5 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_6 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_7 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[3] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_1=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_2=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_3=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_4=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_5=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_6=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_7=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_0 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_1 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_2 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_3 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_4 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_5 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_6 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_7 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[6] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_1=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_2=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_3=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_4=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_5=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_6=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_7=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_0 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_1 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_2 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_3 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_4 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_5 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_6 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_7 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[0] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_1=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_2=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_3=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_4=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_5=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_6=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_7=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_0 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_1 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_2 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_3 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_4 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_5 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_6 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_7 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[5] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_1=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_2=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_3=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_4=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_5=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_6=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_7=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_0 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_1 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_2 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_3 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_4 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_5 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_6 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_7 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[7] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_1=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_2=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_3=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_4=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_5=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_6=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_7=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_0 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_1 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_2 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_3 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_4 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_5 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_6 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_7 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[4] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_1=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_2=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_3=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_4=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_5=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_6=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_7=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_0 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_1 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_2 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_3 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_4 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_5 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_6 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_7 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[2] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_1=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_2=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_3=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_4=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_5=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_6=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_7=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_0 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_1 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_2 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_3 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_4 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_5 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_6 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_7 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[3] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_1=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_2=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_3=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_4=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_5=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_6=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_7=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_0 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_1 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_2 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_3 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_4 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_5 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_6 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_7 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[6] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_1=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_2=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_3=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_4=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_5=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_6=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_7=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_0 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_1 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_2 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_3 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_4 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_5 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_6 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_7 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[0] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_1=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_2=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_3=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_4=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_5=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_6=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_7=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_0 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_1 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_2 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_3 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_4 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_5 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_6 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_7 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[5] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_1=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_2=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_3=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_4=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_5=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_6=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_7=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_0 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_1 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_2 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_3 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_4 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_5 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_6 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_7 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[7] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_1=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_2=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_3=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_4=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_5=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_6=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_7=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_0 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_1 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_2 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_3 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_4 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_5 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_6 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_7 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[4] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_1=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_2=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_3=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_4=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_5=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_6=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_7=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_0 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_1 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_2 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_3 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_4 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_5 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_6 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_7 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[2] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_1=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_2=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_3=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_4=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_5=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_6=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_7=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_0 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_1 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_2 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_3 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_4 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_5 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_6 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_7 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[3] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_1=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_2=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_3=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_4=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_5=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_6=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_7=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_0 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_1 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_2 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_3 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_4 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_5 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_6 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_7 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[6] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_1=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_2=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_3=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_4=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_5=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_6=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_7=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_0 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_1 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_2 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_3 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_4 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_5 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_6 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_7 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[0] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_1=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_2=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_3=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_4=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_5=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_6=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_7=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_0 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_1 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_2 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_3 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_4 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_5 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_6 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_7 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[5] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_1=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_2=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_3=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_4=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_5=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_6=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_7=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_0 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_1 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_2 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_3 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_4 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_5 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_6 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_7 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[7] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_1=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_2=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_3=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_4=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_5=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_6=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_7=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_0 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_1 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_2 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_3 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_4 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_5 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_6 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_7 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[4] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_1=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_2=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_3=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_4=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_5=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_6=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_7=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_0 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_1 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_2 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_3 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_4 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_5 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_6 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_7 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[2] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_1=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_2=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_3=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_4=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_5=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_6=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_7=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_0 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_1 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_2 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_3 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_4 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_5 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_6 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_7 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[3] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_1=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_2=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_3=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_4=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_5=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_6=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_7=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_0 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_1 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_2 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_3 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_4 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_5 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_6 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_7 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[0] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_1=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_2=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_3=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_4=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_5=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_6=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_7=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_0 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_1 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_2 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_3 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_4 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_5 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_6 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_7 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[4] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[4], DdrCtrl_WDATA_0[12], DdrCtrl_WDATA_0[20], 
            DdrCtrl_WDATA_0[28], DdrCtrl_WDATA_0[36], DdrCtrl_WDATA_0[44], 
            DdrCtrl_WDATA_0[52], DdrCtrl_WDATA_0[60], DdrCtrl_WDATA_0[68], 
            DdrCtrl_WDATA_0[76], DdrCtrl_WDATA_0[84], DdrCtrl_WDATA_0[92], 
            DdrCtrl_WDATA_0[100], DdrCtrl_WDATA_0[108], DdrCtrl_WDATA_0[116], 
            DdrCtrl_WDATA_0[124]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[7] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[7], DdrCtrl_WDATA_0[15], DdrCtrl_WDATA_0[23], 
            DdrCtrl_WDATA_0[31], DdrCtrl_WDATA_0[39], DdrCtrl_WDATA_0[47], 
            DdrCtrl_WDATA_0[55], DdrCtrl_WDATA_0[63], DdrCtrl_WDATA_0[71], 
            DdrCtrl_WDATA_0[79], DdrCtrl_WDATA_0[87], DdrCtrl_WDATA_0[95], 
            DdrCtrl_WDATA_0[103], DdrCtrl_WDATA_0[111], DdrCtrl_WDATA_0[119], 
            DdrCtrl_WDATA_0[127]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[6] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[6], DdrCtrl_WDATA_0[14], DdrCtrl_WDATA_0[22], 
            DdrCtrl_WDATA_0[30], DdrCtrl_WDATA_0[38], DdrCtrl_WDATA_0[46], 
            DdrCtrl_WDATA_0[54], DdrCtrl_WDATA_0[62], DdrCtrl_WDATA_0[70], 
            DdrCtrl_WDATA_0[78], DdrCtrl_WDATA_0[86], DdrCtrl_WDATA_0[94], 
            DdrCtrl_WDATA_0[102], DdrCtrl_WDATA_0[110], DdrCtrl_WDATA_0[118], 
            DdrCtrl_WDATA_0[126]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[1] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[1], DdrCtrl_WDATA_0[9], DdrCtrl_WDATA_0[17], 
            DdrCtrl_WDATA_0[25], DdrCtrl_WDATA_0[33], DdrCtrl_WDATA_0[41], 
            DdrCtrl_WDATA_0[49], DdrCtrl_WDATA_0[57], DdrCtrl_WDATA_0[65], 
            DdrCtrl_WDATA_0[73], DdrCtrl_WDATA_0[81], DdrCtrl_WDATA_0[89], 
            DdrCtrl_WDATA_0[97], DdrCtrl_WDATA_0[105], DdrCtrl_WDATA_0[113], 
            DdrCtrl_WDATA_0[121]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[2] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[2], DdrCtrl_WDATA_0[10], DdrCtrl_WDATA_0[18], 
            DdrCtrl_WDATA_0[26], DdrCtrl_WDATA_0[34], DdrCtrl_WDATA_0[42], 
            DdrCtrl_WDATA_0[50], DdrCtrl_WDATA_0[58], DdrCtrl_WDATA_0[66], 
            DdrCtrl_WDATA_0[74], DdrCtrl_WDATA_0[82], DdrCtrl_WDATA_0[90], 
            DdrCtrl_WDATA_0[98], DdrCtrl_WDATA_0[106], DdrCtrl_WDATA_0[114], 
            DdrCtrl_WDATA_0[122]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[0] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[0], DdrCtrl_WDATA_0[8], DdrCtrl_WDATA_0[16], 
            DdrCtrl_WDATA_0[24], DdrCtrl_WDATA_0[32], DdrCtrl_WDATA_0[40], 
            DdrCtrl_WDATA_0[48], DdrCtrl_WDATA_0[56], DdrCtrl_WDATA_0[64], 
            DdrCtrl_WDATA_0[72], DdrCtrl_WDATA_0[80], DdrCtrl_WDATA_0[88], 
            DdrCtrl_WDATA_0[96], DdrCtrl_WDATA_0[104], DdrCtrl_WDATA_0[112], 
            DdrCtrl_WDATA_0[120]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[3] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[3], DdrCtrl_WDATA_0[11], DdrCtrl_WDATA_0[19], 
            DdrCtrl_WDATA_0[27], DdrCtrl_WDATA_0[35], DdrCtrl_WDATA_0[43], 
            DdrCtrl_WDATA_0[51], DdrCtrl_WDATA_0[59], DdrCtrl_WDATA_0[67], 
            DdrCtrl_WDATA_0[75], DdrCtrl_WDATA_0[83], DdrCtrl_WDATA_0[91], 
            DdrCtrl_WDATA_0[99], DdrCtrl_WDATA_0[107], DdrCtrl_WDATA_0[115], 
            DdrCtrl_WDATA_0[123]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[5] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[5], DdrCtrl_WDATA_0[13], DdrCtrl_WDATA_0[21], 
            DdrCtrl_WDATA_0[29], DdrCtrl_WDATA_0[37], DdrCtrl_WDATA_0[45], 
            DdrCtrl_WDATA_0[53], DdrCtrl_WDATA_0[61], DdrCtrl_WDATA_0[69], 
            DdrCtrl_WDATA_0[77], DdrCtrl_WDATA_0[85], DdrCtrl_WDATA_0[93], 
            DdrCtrl_WDATA_0[101], DdrCtrl_WDATA_0[109], DdrCtrl_WDATA_0[117], 
            DdrCtrl_WDATA_0[125]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[4] , 
            \u_axi4_ctrl/rfifo_wdata[12] , \u_axi4_ctrl/rfifo_wdata[20] , 
            \u_axi4_ctrl/rfifo_wdata[28] , \u_axi4_ctrl/rfifo_wdata[36] , 
            \u_axi4_ctrl/rfifo_wdata[44] , \u_axi4_ctrl/rfifo_wdata[52] , 
            \u_axi4_ctrl/rfifo_wdata[60] , \u_axi4_ctrl/rfifo_wdata[68] , 
            \u_axi4_ctrl/rfifo_wdata[76] , \u_axi4_ctrl/rfifo_wdata[84] , 
            \u_axi4_ctrl/rfifo_wdata[92] , \u_axi4_ctrl/rfifo_wdata[100] , 
            \u_axi4_ctrl/rfifo_wdata[108] , \u_axi4_ctrl/rfifo_wdata[116] , 
            \u_axi4_ctrl/rfifo_wdata[124] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[6] , 
            \u_axi4_ctrl/rfifo_wdata[14] , \u_axi4_ctrl/rfifo_wdata[22] , 
            \u_axi4_ctrl/rfifo_wdata[30] , \u_axi4_ctrl/rfifo_wdata[38] , 
            \u_axi4_ctrl/rfifo_wdata[46] , \u_axi4_ctrl/rfifo_wdata[54] , 
            \u_axi4_ctrl/rfifo_wdata[62] , \u_axi4_ctrl/rfifo_wdata[70] , 
            \u_axi4_ctrl/rfifo_wdata[78] , \u_axi4_ctrl/rfifo_wdata[86] , 
            \u_axi4_ctrl/rfifo_wdata[94] , \u_axi4_ctrl/rfifo_wdata[102] , 
            \u_axi4_ctrl/rfifo_wdata[110] , \u_axi4_ctrl/rfifo_wdata[118] , 
            \u_axi4_ctrl/rfifo_wdata[126] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[7] , 
            \u_axi4_ctrl/rfifo_wdata[15] , \u_axi4_ctrl/rfifo_wdata[23] , 
            \u_axi4_ctrl/rfifo_wdata[31] , \u_axi4_ctrl/rfifo_wdata[39] , 
            \u_axi4_ctrl/rfifo_wdata[47] , \u_axi4_ctrl/rfifo_wdata[55] , 
            \u_axi4_ctrl/rfifo_wdata[63] , \u_axi4_ctrl/rfifo_wdata[71] , 
            \u_axi4_ctrl/rfifo_wdata[79] , \u_axi4_ctrl/rfifo_wdata[87] , 
            \u_axi4_ctrl/rfifo_wdata[95] , \u_axi4_ctrl/rfifo_wdata[103] , 
            \u_axi4_ctrl/rfifo_wdata[111] , \u_axi4_ctrl/rfifo_wdata[119] , 
            \u_axi4_ctrl/rfifo_wdata[127] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[2] , 
            \u_axi4_ctrl/rfifo_wdata[10] , \u_axi4_ctrl/rfifo_wdata[18] , 
            \u_axi4_ctrl/rfifo_wdata[26] , \u_axi4_ctrl/rfifo_wdata[34] , 
            \u_axi4_ctrl/rfifo_wdata[42] , \u_axi4_ctrl/rfifo_wdata[50] , 
            \u_axi4_ctrl/rfifo_wdata[58] , \u_axi4_ctrl/rfifo_wdata[66] , 
            \u_axi4_ctrl/rfifo_wdata[74] , \u_axi4_ctrl/rfifo_wdata[82] , 
            \u_axi4_ctrl/rfifo_wdata[90] , \u_axi4_ctrl/rfifo_wdata[98] , 
            \u_axi4_ctrl/rfifo_wdata[106] , \u_axi4_ctrl/rfifo_wdata[114] , 
            \u_axi4_ctrl/rfifo_wdata[122] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[1] , 
            \u_axi4_ctrl/rfifo_wdata[9] , \u_axi4_ctrl/rfifo_wdata[17] , 
            \u_axi4_ctrl/rfifo_wdata[25] , \u_axi4_ctrl/rfifo_wdata[33] , 
            \u_axi4_ctrl/rfifo_wdata[41] , \u_axi4_ctrl/rfifo_wdata[49] , 
            \u_axi4_ctrl/rfifo_wdata[57] , \u_axi4_ctrl/rfifo_wdata[65] , 
            \u_axi4_ctrl/rfifo_wdata[73] , \u_axi4_ctrl/rfifo_wdata[81] , 
            \u_axi4_ctrl/rfifo_wdata[89] , \u_axi4_ctrl/rfifo_wdata[97] , 
            \u_axi4_ctrl/rfifo_wdata[105] , \u_axi4_ctrl/rfifo_wdata[113] , 
            \u_axi4_ctrl/rfifo_wdata[121] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[0] , 
            \u_axi4_ctrl/rfifo_wdata[8] , \u_axi4_ctrl/rfifo_wdata[16] , 
            \u_axi4_ctrl/rfifo_wdata[24] , \u_axi4_ctrl/rfifo_wdata[32] , 
            \u_axi4_ctrl/rfifo_wdata[40] , \u_axi4_ctrl/rfifo_wdata[48] , 
            \u_axi4_ctrl/rfifo_wdata[56] , \u_axi4_ctrl/rfifo_wdata[64] , 
            \u_axi4_ctrl/rfifo_wdata[72] , \u_axi4_ctrl/rfifo_wdata[80] , 
            \u_axi4_ctrl/rfifo_wdata[88] , \u_axi4_ctrl/rfifo_wdata[96] , 
            \u_axi4_ctrl/rfifo_wdata[104] , \u_axi4_ctrl/rfifo_wdata[112] , 
            \u_axi4_ctrl/rfifo_wdata[120] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[3] , 
            \u_axi4_ctrl/rfifo_wdata[11] , \u_axi4_ctrl/rfifo_wdata[19] , 
            \u_axi4_ctrl/rfifo_wdata[27] , \u_axi4_ctrl/rfifo_wdata[35] , 
            \u_axi4_ctrl/rfifo_wdata[43] , \u_axi4_ctrl/rfifo_wdata[51] , 
            \u_axi4_ctrl/rfifo_wdata[59] , \u_axi4_ctrl/rfifo_wdata[67] , 
            \u_axi4_ctrl/rfifo_wdata[75] , \u_axi4_ctrl/rfifo_wdata[83] , 
            \u_axi4_ctrl/rfifo_wdata[91] , \u_axi4_ctrl/rfifo_wdata[99] , 
            \u_axi4_ctrl/rfifo_wdata[107] , \u_axi4_ctrl/rfifo_wdata[115] , 
            \u_axi4_ctrl/rfifo_wdata[123] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[5] , 
            \u_axi4_ctrl/rfifo_wdata[13] , \u_axi4_ctrl/rfifo_wdata[21] , 
            \u_axi4_ctrl/rfifo_wdata[29] , \u_axi4_ctrl/rfifo_wdata[37] , 
            \u_axi4_ctrl/rfifo_wdata[45] , \u_axi4_ctrl/rfifo_wdata[53] , 
            \u_axi4_ctrl/rfifo_wdata[61] , \u_axi4_ctrl/rfifo_wdata[69] , 
            \u_axi4_ctrl/rfifo_wdata[77] , \u_axi4_ctrl/rfifo_wdata[85] , 
            \u_axi4_ctrl/rfifo_wdata[93] , \u_axi4_ctrl/rfifo_wdata[101] , 
            \u_axi4_ctrl/rfifo_wdata[109] , \u_axi4_ctrl/rfifo_wdata[117] , 
            \u_axi4_ctrl/rfifo_wdata[125] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[8] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=50250a83 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[9] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=b3ca6a06 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=f7222e73 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[10] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=e72ac1a0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=b985acac */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=7af58ba3 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=451f771f */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=19baebb3 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=b9119f89 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=5b8fe925 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12  (.WCLK(\tx_slowclk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n661 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=a4bb9c7d */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity/work_dbg/debug_top.v(410)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .READ_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, n1175, n1176, n1178, n1180, 
            n1182, n1199, n1201, n1203, n1205, n1207, n1209, n1731}), 
            .B({10'b0000000000, \u_scaler_gray/tdata01[7] , \u_scaler_gray/tdata01[6] , 
            \u_scaler_gray/tdata01[5] , \u_scaler_gray/tdata01[4] , \u_scaler_gray/tdata01[3] , 
            \u_scaler_gray/tdata01[2] , \u_scaler_gray/tdata01[1] , \u_scaler_gray/tdata01[0] }), 
            .O({Open_0, Open_1, Open_2, Open_3, Open_4, Open_5, 
            Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, Open_12, 
            Open_13, Open_14, Open_15, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[19] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[18] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[17] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[16] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[15] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[14] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[13] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[12] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[11] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[10] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[9] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[8] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[7] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[6] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[5] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[4] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[3] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[2] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[1] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(33)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, n1154, n1155, n1157, n1159, 
            n1161, n1163, n1165, n1167, n1169, n1171, n1173, n1733}), 
            .B({10'b0000000000, \u_scaler_gray/tdata10[7] , \u_scaler_gray/tdata10[6] , 
            \u_scaler_gray/tdata10[5] , \u_scaler_gray/tdata10[4] , \u_scaler_gray/tdata10[3] , 
            \u_scaler_gray/tdata10[2] , \u_scaler_gray/tdata10[1] , \u_scaler_gray/tdata10[0] }), 
            .O({Open_16, Open_17, Open_18, Open_19, Open_20, Open_21, 
            Open_22, Open_23, Open_24, Open_25, Open_26, Open_27, 
            Open_28, Open_29, Open_30, Open_31, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[19] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[18] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[17] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[16] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[15] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[14] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[13] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[12] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[11] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[10] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[9] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[8] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[7] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[6] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[5] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[4] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[3] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[2] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[1] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(34)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b0), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] }), 
            .B({6'b000000, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0] }), 
            .O({Open_32, Open_33, Open_34, Open_35, Open_36, Open_37, 
            Open_38, Open_39, Open_40, Open_41, Open_42, Open_43, 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[23] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[22] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[21] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[20] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[19] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[18] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[17] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[16] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[15] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[14] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[13] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[12] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[11] , 
            Open_44, Open_45, Open_46, Open_47, Open_48, Open_49, 
            Open_50, Open_51, Open_52, Open_53, Open_54})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b0, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b0, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(50)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .A_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTA_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b0), .RSTA(1'b0), .CEB(1'b1), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] }), 
            .B({6'b000000, \u_scaler_gray/u1_bilinear_gray/srcy_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[10] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[8] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[7] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[6] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[5] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[4] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[3] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[2] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[1] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[0] }), .O({Open_55, 
            Open_56, Open_57, Open_58, Open_59, Open_60, Open_61, 
            Open_62, Open_63, Open_64, Open_65, Open_66, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[23] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[22] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[21] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[20] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[19] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[18] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[17] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[16] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[15] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[14] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[13] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[12] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[11] , 
            Open_67, Open_68, Open_69, Open_70, Open_71, Open_72, 
            Open_73, Open_74, Open_75, Open_76, Open_77})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b0, B_REG=1'b1, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b0, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b1, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(52)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .A_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .B_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTA_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTB_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b0), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({18'b000001001100110011}), .B({2'b00, \u_scaler_gray/desty[15] , 
            \u_scaler_gray/desty[14] , \u_scaler_gray/desty[13] , \u_scaler_gray/desty[12] , 
            \u_scaler_gray/desty[11] , \u_scaler_gray/desty[10] , \u_scaler_gray/desty[9] , 
            \u_scaler_gray/desty[8] , \u_scaler_gray/desty[7] , \u_scaler_gray/desty[6] , 
            \u_scaler_gray/desty[5] , \u_scaler_gray/desty[4] , \u_scaler_gray/desty[3] , 
            \u_scaler_gray/desty[2] , \u_scaler_gray/desty[1] , \u_scaler_gray/desty[0] }), 
            .O({Open_78, Open_79, Open_80, Open_81, Open_82, Open_83, 
            Open_84, Open_85, \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[27] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[26] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[25] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[24] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[23] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[22] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[21] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[20] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[19] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[18] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[17] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[16] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[15] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[14] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[13] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[12] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[11] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[10] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[9] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[8] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[7] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[6] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[5] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[4] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[3] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[2] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[1] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b0, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b0, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(55)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .A_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTA_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, n1211, n1212, n1214, n1216, 
            n1218, n1220, n1222, n1224, n1226, n1228, n1230, n1688}), 
            .B({10'b0000000000, \u_scaler_gray/tdata00[7] , \u_scaler_gray/tdata00[6] , 
            \u_scaler_gray/tdata00[5] , \u_scaler_gray/tdata00[4] , \u_scaler_gray/tdata00[3] , 
            \u_scaler_gray/tdata00[2] , \u_scaler_gray/tdata00[1] , \u_scaler_gray/tdata00[0] }), 
            .O({Open_86, Open_87, Open_88, Open_89, Open_90, Open_91, 
            Open_92, Open_93, Open_94, Open_95, Open_96, Open_97, 
            Open_98, Open_99, Open_100, Open_101, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[19] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[18] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[17] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[16] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[15] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[14] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[13] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[12] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[11] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[10] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[9] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[8] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[7] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[6] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[5] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[4] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[3] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[2] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[1] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(32)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b1), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, \u_scaler_gray/u1_bilinear_gray/srcx_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/srcx_fix[10] , \u_scaler_gray/u1_bilinear_gray/srcx_fix[9] , 
            9'b000000000}), .B({6'b000000, \u_scaler_gray/u1_bilinear_gray/srcy_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[10] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[8] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[7] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[6] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[5] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[4] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[3] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[2] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[1] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[0] }), .O({Open_102, 
            Open_103, Open_104, Open_105, Open_106, Open_107, Open_108, 
            Open_109, Open_110, Open_111, Open_112, Open_113, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[23] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[22] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[21] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[20] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[19] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[18] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[17] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[16] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[15] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[14] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[13] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[12] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[11] , 
            Open_114, Open_115, Open_116, Open_117, Open_118, Open_119, 
            Open_120, Open_121, Open_122, Open_123, Open_124})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b1, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b1, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(53)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .B_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTB_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, \u_scaler_gray/u1_bilinear_gray/srcx_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/srcx_fix[10] , \u_scaler_gray/u1_bilinear_gray/srcx_fix[9] , 
            9'b000000000}), .B({6'b000000, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0] }), 
            .O({Open_125, Open_126, Open_127, Open_128, Open_129, 
            Open_130, Open_131, Open_132, Open_133, Open_134, Open_135, 
            Open_136, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[23] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[22] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[21] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[20] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[19] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[18] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[17] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[16] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[15] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[14] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[13] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[12] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[11] , 
            Open_137, Open_138, Open_139, Open_140, Open_141, Open_142, 
            Open_143, Open_144, Open_145, Open_146, Open_147})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(51)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, n1133, n1134, n1136, n1138, 
            n1140, n1142, n1144, n1146, n1148, n1150, n1152, n1735}), 
            .B({10'b0000000000, \u_scaler_gray/tdata11[7] , \u_scaler_gray/tdata11[6] , 
            \u_scaler_gray/tdata11[5] , \u_scaler_gray/tdata11[4] , \u_scaler_gray/tdata11[3] , 
            \u_scaler_gray/tdata11[2] , \u_scaler_gray/tdata11[1] , \u_scaler_gray/tdata11[0] }), 
            .O({Open_148, Open_149, Open_150, Open_151, Open_152, 
            Open_153, Open_154, Open_155, Open_156, Open_157, Open_158, 
            Open_159, Open_160, Open_161, Open_162, Open_163, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[19] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[18] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[17] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[16] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[15] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[14] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[13] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[12] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[11] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[10] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[9] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[8] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[7] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[6] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[5] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[4] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[3] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[2] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[1] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__15142 (.I0(\u_axi4_ctrl/wdata_cnt_dly[4] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[5] ), 
            .I2(n10069), .O(n10070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15142.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15143 (.I0(\u_axi4_ctrl/wdata_cnt_dly[2] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[3] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[4] ), .I3(\u_axi4_ctrl/wdata_cnt_dly[5] ), 
            .O(n10071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15143.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15144 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(n10071), .O(n10072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15144.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15145 (.I0(n10072), .I1(n10070), .I2(DdrCtrl_WREADY_0), 
            .I3(\u_axi4_ctrl/wdata_cnt_dly[6] ), .O(n10073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__15145.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__15146 (.I0(\u_axi4_ctrl/state[2] ), .I1(\u_axi4_ctrl/state[1] ), 
            .O(DdrCtrl_BREADY_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15146.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15147 (.I0(\u_axi4_ctrl/state[0] ), .I1(DdrCtrl_BREADY_0), 
            .O(DdrCtrl_WVALID_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15147.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15148 (.I0(\u_axi4_ctrl/wdata_cnt_dly[7] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[8] ), 
            .I2(n10073), .I3(DdrCtrl_WVALID_0), .O(DdrCtrl_WLAST_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15148.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15149 (.I0(\u_axi4_ctrl/state[1] ), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(\u_axi4_ctrl/state[2] ), .O(DdrCtrl_RREADY_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15149.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15150 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), .O(n10074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h45fe */ ;
    defparam LUT__15150.LUTMASK = 16'h45fe;
    EFX_LUT4 LUT__15151 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), .O(n10075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfd3f */ ;
    defparam LUT__15151.LUTMASK = 16'hfd3f;
    EFX_LUT4 LUT__15152 (.I0(n10074), .I1(n10075), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk ), 
            .O(cmos_sclk)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__15152.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__15153 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .O(n10076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15153.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15154 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I1(n10076), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I3(n10074), .O(cmos_sdat_OE)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bff */ ;
    defparam LUT__15154.LUTMASK = 16'h0bff;
    EFX_LUT4 LUT__15155 (.I0(\PowerOnResetCnt[4] ), .I1(\PowerOnResetCnt[5] ), 
            .I2(\PowerOnResetCnt[6] ), .I3(\PowerOnResetCnt[7] ), .O(n10077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15155.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15156 (.I0(\PowerOnResetCnt[0] ), .I1(\PowerOnResetCnt[1] ), 
            .I2(\PowerOnResetCnt[2] ), .I3(\PowerOnResetCnt[3] ), .O(n10078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15156.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15157 (.I0(n10077), .I1(n10078), .O(\reduce_nand_9/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15157.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15158 (.I0(\r_hdmi_tx0_o[5] ), .I1(\w_hdmi_txd0[0] ), 
            .I2(rc_hdmi_tx), .O(n592_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15158.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15159 (.I0(\r_hdmi_tx1_o[5] ), .I1(\w_hdmi_txd1[0] ), 
            .I2(rc_hdmi_tx), .O(n603_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15159.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15160 (.I0(\r_hdmi_tx2_o[5] ), .I1(\w_hdmi_txd2[0] ), 
            .I2(rc_hdmi_tx), .O(n614_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15160.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15161 (.I0(PllLocked[1]), .I1(PllLocked[0]), .O(n9_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15161.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15162 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] ), .O(n10079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15162.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15163 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] ), .O(n10080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15163.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15164 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] ), .O(n10081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15164.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15165 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] ), .O(n10082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15165.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15166 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] ), .O(n10083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15166.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15167 (.I0(n10080), .I1(n10081), .I2(n10082), .I3(n10083), 
            .O(n10084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15167.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15168 (.I0(n10079), .I1(n10084), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__15168.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__15169 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/equal_21/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__15169.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__15170 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__15170.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__15171 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__15171.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__15172 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3] ), .O(n10085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15172.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15173 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] ), .I2(n10085), 
            .O(n10086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15173.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15174 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] ), 
            .I1(n10086), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] ), .O(n10087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__15174.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__15175 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), .O(n10088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15175.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15176 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), 
            .I1(n10087), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), 
            .I3(n10088), .O(n10089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__15176.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__15177 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11] ), .O(n10090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__15177.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__15178 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14] ), 
            .O(n10091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15178.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15179 (.I0(n10090), .I1(n10091), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16] ), .O(n10092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__15179.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__15180 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11] ), .O(n10093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15180.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15181 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15] ), .I2(n10093), 
            .O(n10094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15181.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15182 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19] ), 
            .O(n10095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15182.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15183 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4] ), .O(n10096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15183.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15184 (.I0(n10092), .I1(n10094), .I2(n10095), .I3(n10096), 
            .O(n10097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15184.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15185 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15] ), .I2(n10097), 
            .O(n10098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15185.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15186 (.I0(n10089), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13] ), 
            .I2(n10098), .O(n10099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15186.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15187 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] ), 
            .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15187.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15188 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3] ), .O(n10100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15188.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15189 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I3(n10100), .O(n10101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__15189.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__15190 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .O(n10102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15190.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15191 (.I0(n10102), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), .O(n10103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15191.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15192 (.I0(n10103), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .O(n10104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__15192.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__15193 (.I0(n10101), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .I3(n10104), 
            .O(n10105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__15193.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__15194 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[6] ), 
            .I2(\i2c_config_index[7] ), .O(n10106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15194.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15195 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[3] ), 
            .I2(n10106), .O(n10107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__15195.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__15196 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I3(n10107), .O(n10108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15196.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15197 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .O(n10109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__15197.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__15198 (.I0(n10109), .I1(n10100), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .O(n10110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15198.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15199 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), 
            .O(n10111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__15199.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__15200 (.I0(n10097), .I1(n10108), .I2(n10110), .I3(n10111), 
            .O(n10112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__15200.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__15201 (.I0(n10105), .I1(n10112), .O(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__15201.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__15202 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3] ), .O(n10113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15202.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15203 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4] ), 
            .I1(n10113), .O(n10114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15203.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15204 (.I0(n10114), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] ), 
            .O(n10115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15204.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15205 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] ), 
            .I1(n10115), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] ), .O(n10116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__15205.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__15206 (.I0(n10116), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] ), 
            .O(n10117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__15206.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__15207 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] ), .O(n10118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15207.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15208 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), .I2(n10115), 
            .I3(n10118), .O(n10119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15208.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15209 (.I0(n10119), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), 
            .O(n10120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15209.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15210 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13] ), 
            .I1(n10098), .O(n10121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15210.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15211 (.I0(n10117), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), 
            .I2(n10120), .I3(n10121), .O(\u_i2c_timing_ctrl_16reg_16bit/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__15211.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__15212 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] ), .I2(n10121), 
            .I3(n10118), .O(n10122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15212.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15213 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), .O(n10123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15213.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15214 (.I0(n10114), .I1(n10122), .I2(n10123), .O(\u_i2c_timing_ctrl_16reg_16bit/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15214.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15215 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), 
            .I3(n10086), .O(n10124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15215.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15216 (.I0(n10122), .I1(n10124), .O(\u_i2c_timing_ctrl_16reg_16bit/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15216.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15217 (.I0(\i2c_config_index[0] ), .I1(n10107), .O(\u_i2c_timing_ctrl_16reg_16bit/n205 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15217.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15218 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), .O(n10125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15218.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15219 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack ), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .O(n10126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__15219.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__15220 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .I2(n10125), 
            .I3(n10126), .O(\u_i2c_timing_ctrl_16reg_16bit/n846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15220.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15221 (.I0(n10100), .I1(n10076), .I2(n10102), .O(n10127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15221.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15222 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I1(n10102), .O(n10128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15222.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15223 (.I0(n10125), .I1(n10101), .I2(n10128), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .O(n10129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbaf0 */ ;
    defparam LUT__15223.LUTMASK = 16'hbaf0;
    EFX_LUT4 LUT__15224 (.I0(n10127), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I2(n10129), .O(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__15224.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__15225 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), 
            .O(n10130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15225.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15226 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[0] ), .O(n10131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ffa */ ;
    defparam LUT__15226.LUTMASK = 16'h3ffa;
    EFX_LUT4 LUT__15227 (.I0(n10131), .I1(n10106), .O(n10132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15227.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15228 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[4] ), 
            .O(n10133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15228.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15229 (.I0(n10130), .I1(n10132), .I2(n10133), .O(n10134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15229.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15230 (.I0(n10097), .I1(n10134), .I2(n10128), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .O(n10135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ff8 */ ;
    defparam LUT__15230.LUTMASK = 16'h0ff8;
    EFX_LUT4 LUT__15231 (.I0(n10130), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .O(n10136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__15231.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__15232 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I1(n10102), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I3(n10100), .O(n10137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h570f */ ;
    defparam LUT__15232.LUTMASK = 16'h570f;
    EFX_LUT4 LUT__15233 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I3(n10102), .O(n10138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbaf0 */ ;
    defparam LUT__15233.LUTMASK = 16'hbaf0;
    EFX_LUT4 LUT__15234 (.I0(n10137), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I2(n10138), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .O(n10139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__15234.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__15235 (.I0(n10136), .I1(n10135), .I2(n10139), .O(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8 */ ;
    defparam LUT__15235.LUTMASK = 16'hf8f8;
    EFX_LUT4 LUT__15236 (.I0(n10097), .I1(n10134), .O(n10140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15236.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15237 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I1(n10130), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I3(n10128), .O(n10141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0230 */ ;
    defparam LUT__15237.LUTMASK = 16'h0230;
    EFX_LUT4 LUT__15238 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I1(n10140), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I3(n10141), .O(n10142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__15238.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__15239 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I1(n10137), .O(n10143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15239.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15240 (.I0(n10143), .I1(n10104), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .I3(n10142), .O(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h444f */ ;
    defparam LUT__15240.LUTMASK = 16'h444f;
    EFX_LUT4 LUT__15241 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__15241.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__15242 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), .O(n10145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15242.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15243 (.I0(n10125), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I2(n10102), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5780 */ ;
    defparam LUT__15243.LUTMASK = 16'h5780;
    EFX_LUT4 LUT__15244 (.I0(n10144), .I1(n10145), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), .O(n10146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3fa */ ;
    defparam LUT__15244.LUTMASK = 16'hc3fa;
    EFX_LUT4 LUT__15245 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I1(n10146), .O(\u_i2c_timing_ctrl_16reg_16bit/n500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15245.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15246 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), .O(n10147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h32f3 */ ;
    defparam LUT__15246.LUTMASK = 16'h32f3;
    EFX_LUT4 LUT__15247 (.I0(n10147), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .O(ceg_net552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15247.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15248 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), .O(n10148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1004 */ ;
    defparam LUT__15248.LUTMASK = 16'h1004;
    EFX_LUT4 LUT__15249 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[2] ), .O(n10149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7fe */ ;
    defparam LUT__15249.LUTMASK = 16'he7fe;
    EFX_LUT4 LUT__15250 (.I0(\i2c_config_index[1] ), .I1(n10149), .I2(n10106), 
            .O(n10150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15250.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15251 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[4] ), .I3(n10106), .O(n10151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15251.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15252 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .I2(n10151), .O(n10152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15252.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15253 (.I0(n10152), .I1(n10150), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .O(n10153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15253.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15254 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(n10152), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), .O(n10154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__15254.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__15255 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[2] ), .O(n10155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hdcab */ ;
    defparam LUT__15255.LUTMASK = 16'hdcab;
    EFX_LUT4 LUT__15256 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[4] ), .O(n10156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__15256.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__15257 (.I0(\i2c_config_index[0] ), .I1(n10156), .I2(\i2c_config_index[2] ), 
            .O(n10157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15257.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15258 (.I0(n10155), .I1(\i2c_config_index[1] ), .I2(n10157), 
            .I3(n10106), .O(n10158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__15258.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__15259 (.I0(n10158), .I1(n10154), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .O(n10159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__15259.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__15260 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(n10153), .I2(n10159), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77 */ ;
    defparam LUT__15260.LUTMASK = 16'h0f77;
    EFX_LUT4 LUT__15261 (.I0(n10148), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0] ), 
            .I2(n10160), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h440f */ ;
    defparam LUT__15261.LUTMASK = 16'h440f;
    EFX_LUT4 LUT__15262 (.I0(n10142), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .O(n10161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15262.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15263 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .O(n10162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15263.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15264 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), .I2(n10162), 
            .O(n10163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__15264.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__15265 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .I1(n10163), .I2(n10161), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), 
            .O(ceg_net664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__15265.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__15266 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), .O(n10164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15266.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15267 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(n10162), .I2(n10164), .O(n10165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15267.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15268 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), .O(n10166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15268.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15269 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I3(n10166), .O(n10167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15269.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15270 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack5 ), .I1(cmos_sdat_IN), 
            .I2(n10165), .I3(n10167), .O(\u_i2c_timing_ctrl_16reg_16bit/n567 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcfa */ ;
    defparam LUT__15270.LUTMASK = 16'hfcfa;
    EFX_LUT4 LUT__15271 (.I0(n10105), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I2(n10162), .O(n10168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15271.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15272 (.I0(n10164), .I1(cmos_sdat_IN), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack4 ), 
            .I3(n10168), .O(n10169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__15272.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__15273 (.I0(n10163), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack4 ), 
            .I2(n10164), .I3(n10169), .O(\u_i2c_timing_ctrl_16reg_16bit/n570 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ff */ ;
    defparam LUT__15273.LUTMASK = 16'he0ff;
    EFX_LUT4 LUT__15274 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .I3(n10166), .O(n10170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400 */ ;
    defparam LUT__15274.LUTMASK = 16'h1400;
    EFX_LUT4 LUT__15275 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack3 ), .I1(cmos_sdat_IN), 
            .I2(n10165), .I3(n10170), .O(\u_i2c_timing_ctrl_16reg_16bit/n573 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcfa */ ;
    defparam LUT__15275.LUTMASK = 16'hfcfa;
    EFX_LUT4 LUT__15276 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), .O(n10171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15276.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15277 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .I3(n10171), .O(n10172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400 */ ;
    defparam LUT__15277.LUTMASK = 16'h1400;
    EFX_LUT4 LUT__15278 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack2 ), .I1(cmos_sdat_IN), 
            .I2(n10165), .I3(n10172), .O(\u_i2c_timing_ctrl_16reg_16bit/n576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcfa */ ;
    defparam LUT__15278.LUTMASK = 16'hfcfa;
    EFX_LUT4 LUT__15279 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I3(n10166), .O(n10173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100 */ ;
    defparam LUT__15279.LUTMASK = 16'h4100;
    EFX_LUT4 LUT__15280 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack1 ), .I1(cmos_sdat_IN), 
            .I2(n10165), .I3(n10173), .O(\u_i2c_timing_ctrl_16reg_16bit/n579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcfa */ ;
    defparam LUT__15280.LUTMASK = 16'hfcfa;
    EFX_LUT4 LUT__15281 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack4 ), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack3 ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack2 ), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack1 ), 
            .O(n10174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15281.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15282 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack5 ), .I2(n10174), 
            .O(n10175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15282.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15283 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .I1(n10139), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I3(n10144), .O(n10176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__15283.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__15284 (.I0(n10175), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack ), 
            .I2(n10165), .I3(n10176), .O(\u_i2c_timing_ctrl_16reg_16bit/n581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf5fc */ ;
    defparam LUT__15284.LUTMASK = 16'hf5fc;
    EFX_LUT4 LUT__15285 (.I0(n10092), .I1(n10095), .O(\u_i2c_timing_ctrl_16reg_16bit/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15285.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15286 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .O(n10177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__15286.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__15287 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I3(n10177), .O(n10178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__15287.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__15288 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .O(n10179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__15288.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__15289 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I3(n10179), .O(n10180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__15289.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__15290 (.I0(n10180), .I1(n10178), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] ), 
            .O(n10181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15290.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15291 (.I0(n10181), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .O(n10182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15291.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15292 (.I0(n10145), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), .I3(n10182), 
            .O(n10183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__15292.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__15293 (.I0(cmos_sdat_OUT), .I1(n10166), .O(n10184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15293.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15294 (.I0(n10184), .I1(n10162), .I2(n10181), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h15cf */ ;
    defparam LUT__15294.LUTMASK = 16'h15cf;
    EFX_LUT4 LUT__15295 (.I0(n10181), .I1(cmos_sdat_OUT), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), .O(n10186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__15295.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__15296 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] ), 
            .O(n10187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15296.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15297 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3] ), 
            .I1(n10187), .O(n10188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15297.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15298 (.I0(n10188), .I1(n10182), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .O(n10189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__15298.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__15299 (.I0(cmos_sdat_OUT), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .O(n10190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h57c5 */ ;
    defparam LUT__15299.LUTMASK = 16'h57c5;
    EFX_LUT4 LUT__15300 (.I0(n10189), .I1(n10186), .I2(n10190), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__15300.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__15301 (.I0(n10183), .I1(n10185), .I2(n10191), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__15301.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__15302 (.I0(n10112), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I2(n10162), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), 
            .O(ceg_net632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7d00 */ ;
    defparam LUT__15302.LUTMASK = 16'h7d00;
    EFX_LUT4 LUT__15303 (.I0(n228), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15303.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15304 (.I0(n3348), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15304.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15305 (.I0(n3346), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15305.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15306 (.I0(n3341), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15306.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15307 (.I0(n3337), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15307.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15308 (.I0(n3335), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15308.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15309 (.I0(n3333), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15309.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15310 (.I0(n3331), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15310.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15311 (.I0(n3329), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15311.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15312 (.I0(n3323), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15312.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15313 (.I0(n3321), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15313.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15314 (.I0(n3319), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15314.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15315 (.I0(n3317), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15315.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15316 (.I0(n3306), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15316.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15317 (.I0(n3305), .I1(n10099), .O(\u_i2c_timing_ctrl_16reg_16bit/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15317.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15318 (.I0(n231), .I1(n10107), .O(\u_i2c_timing_ctrl_16reg_16bit/n204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15318.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15319 (.I0(n3303), .I1(n10107), .O(\u_i2c_timing_ctrl_16reg_16bit/n203 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15319.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15320 (.I0(n3301), .I1(n10107), .O(\u_i2c_timing_ctrl_16reg_16bit/n202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__15320.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__15321 (.I0(n3299), .I1(n10107), .O(\u_i2c_timing_ctrl_16reg_16bit/n201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__15321.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__15322 (.I0(n3297), .I1(n10107), .O(\u_i2c_timing_ctrl_16reg_16bit/n200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15322.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15323 (.I0(n3295), .I1(n10107), .O(\u_i2c_timing_ctrl_16reg_16bit/n199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15323.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15324 (.I0(n3294), .I1(n10107), .O(\u_i2c_timing_ctrl_16reg_16bit/n198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15324.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15325 (.I0(n10146), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .O(\u_i2c_timing_ctrl_16reg_16bit/n499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__15325.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__15326 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .I2(n10146), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] ), .O(\u_i2c_timing_ctrl_16reg_16bit/n498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__15326.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__15327 (.I0(n10146), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3] ), 
            .I2(n10187), .O(\u_i2c_timing_ctrl_16reg_16bit/n497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__15327.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__15328 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), .O(n10192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__15328.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__15329 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[4] ), .O(n10193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4ccf */ ;
    defparam LUT__15329.LUTMASK = 16'h4ccf;
    EFX_LUT4 LUT__15330 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[0] ), .O(n10194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc17 */ ;
    defparam LUT__15330.LUTMASK = 16'hfc17;
    EFX_LUT4 LUT__15331 (.I0(n10194), .I1(\i2c_config_index[4] ), .I2(\i2c_config_index[3] ), 
            .I3(n10193), .O(n10195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heee0 */ ;
    defparam LUT__15331.LUTMASK = 16'heee0;
    EFX_LUT4 LUT__15332 (.I0(n10195), .I1(n10106), .O(n10196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15332.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15333 (.I0(n10196), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] ), 
            .I2(n10171), .O(n10197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15333.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15334 (.I0(n10197), .I1(n10145), .I2(n10192), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] ), 
            .O(n10198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__15334.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__15335 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[4] ), .O(n10199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb4f */ ;
    defparam LUT__15335.LUTMASK = 16'hfb4f;
    EFX_LUT4 LUT__15336 (.I0(n10199), .I1(n10106), .I2(\i2c_config_index[2] ), 
            .O(n10200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15336.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15337 (.I0(n10196), .I1(n10200), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .O(n10201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15337.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15338 (.I0(\i2c_config_index[3] ), .I1(n10194), .I2(\i2c_config_index[2] ), 
            .I3(n10107), .O(n10202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__15338.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__15339 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] ), .I2(n10202), 
            .I3(n10161), .O(n10203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__15339.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__15340 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I1(n10201), .I2(n10203), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077 */ ;
    defparam LUT__15340.LUTMASK = 16'hf077;
    EFX_LUT4 LUT__15341 (.I0(n10204), .I1(n10198), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15341.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15342 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[2] ), .O(n10205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1700 */ ;
    defparam LUT__15342.LUTMASK = 16'h1700;
    EFX_LUT4 LUT__15343 (.I0(n10199), .I1(n10205), .I2(\i2c_config_index[0] ), 
            .I3(n10106), .O(n10206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1c00 */ ;
    defparam LUT__15343.LUTMASK = 16'h1c00;
    EFX_LUT4 LUT__15344 (.I0(n10206), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] ), 
            .I2(n10171), .O(n10207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15344.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15345 (.I0(n10207), .I1(n10145), .I2(n10192), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] ), 
            .O(n10208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__15345.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__15346 (.I0(\i2c_config_index[4] ), .I1(n10132), .I2(n10206), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), .O(n10209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__15346.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__15347 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[0] ), 
            .O(n10210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15347.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15348 (.I0(\i2c_config_index[2] ), .I1(n10210), .O(n10211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15348.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15349 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[2] ), .O(n10212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3001 */ ;
    defparam LUT__15349.LUTMASK = 16'h3001;
    EFX_LUT4 LUT__15350 (.I0(n10212), .I1(n10211), .I2(\i2c_config_index[1] ), 
            .I3(n10106), .O(n10213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__15350.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__15351 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] ), .I2(n10213), 
            .I3(n10161), .O(n10214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__15351.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__15352 (.I0(n10209), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I2(n10214), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__15352.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__15353 (.I0(n10215), .I1(n10208), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15353.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15354 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), .I2(n10171), 
            .O(n10216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15354.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15355 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[3] ), .O(n10217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3207 */ ;
    defparam LUT__15355.LUTMASK = 16'h3207;
    EFX_LUT4 LUT__15356 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[4] ), .I3(n10210), .O(n10218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc700 */ ;
    defparam LUT__15356.LUTMASK = 16'hc700;
    EFX_LUT4 LUT__15357 (.I0(\i2c_config_index[2] ), .I1(n10217), .I2(n10218), 
            .I3(n10106), .O(n10219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__15357.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__15358 (.I0(n10216), .I1(n10219), .I2(n10148), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3] ), 
            .O(n10220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__15358.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__15359 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .O(n10221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15359.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15360 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[3] ), .O(n10222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa3f */ ;
    defparam LUT__15360.LUTMASK = 16'hfa3f;
    EFX_LUT4 LUT__15361 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[3] ), .O(n10223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15361.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15362 (.I0(\i2c_config_index[4] ), .I1(n10223), .I2(\i2c_config_index[0] ), 
            .O(n10224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15362.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15363 (.I0(n10222), .I1(\i2c_config_index[1] ), .I2(n10224), 
            .I3(n10106), .O(n10225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__15363.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__15364 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3] ), .I2(n10225), 
            .I3(n10161), .O(n10226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__15364.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__15365 (.I0(n10221), .I1(n10219), .I2(n10226), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077 */ ;
    defparam LUT__15365.LUTMASK = 16'hf077;
    EFX_LUT4 LUT__15366 (.I0(n10227), .I1(n10220), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15366.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15367 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[1] ), .O(n10228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe3f */ ;
    defparam LUT__15367.LUTMASK = 16'hfe3f;
    EFX_LUT4 LUT__15368 (.I0(n10228), .I1(\i2c_config_index[2] ), .I2(n10107), 
            .O(n10229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__15368.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__15369 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(n10229), .O(n10230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15369.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15370 (.I0(n10230), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .O(n10231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__15370.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__15371 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[4] ), .O(n10232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ff2 */ ;
    defparam LUT__15371.LUTMASK = 16'h3ff2;
    EFX_LUT4 LUT__15372 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[4] ), .O(n10233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd08c */ ;
    defparam LUT__15372.LUTMASK = 16'hd08c;
    EFX_LUT4 LUT__15373 (.I0(n10232), .I1(n10233), .I2(\i2c_config_index[3] ), 
            .I3(n10106), .O(n10234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1c00 */ ;
    defparam LUT__15373.LUTMASK = 16'h1c00;
    EFX_LUT4 LUT__15374 (.I0(n10205), .I1(\i2c_config_index[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I3(n10234), .O(n10235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15374.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15375 (.I0(n10235), .I1(n10231), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), .O(n10236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccc5 */ ;
    defparam LUT__15375.LUTMASK = 16'hccc5;
    EFX_LUT4 LUT__15376 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[3] ), .O(n10237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe35 */ ;
    defparam LUT__15376.LUTMASK = 16'hfe35;
    EFX_LUT4 LUT__15377 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[4] ), 
            .I2(n10131), .I3(n10237), .O(n10238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc45 */ ;
    defparam LUT__15377.LUTMASK = 16'hfc45;
    EFX_LUT4 LUT__15378 (.I0(n10238), .I1(n10106), .I2(n10230), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__15378.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__15379 (.I0(n10239), .I1(n10236), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), .O(n10240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hccca */ ;
    defparam LUT__15379.LUTMASK = 16'hccca;
    EFX_LUT4 LUT__15380 (.I0(n10234), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4] ), 
            .I2(n10171), .I3(n10145), .O(n10241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__15380.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__15381 (.I0(n10241), .I1(n10192), .I2(n10240), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hab0f */ ;
    defparam LUT__15381.LUTMASK = 16'hab0f;
    EFX_LUT4 LUT__15382 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[3] ), .O(n10242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe4f */ ;
    defparam LUT__15382.LUTMASK = 16'hfe4f;
    EFX_LUT4 LUT__15383 (.I0(n10242), .I1(n10133), .I2(\i2c_config_index[2] ), 
            .I3(n10106), .O(n10243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__15383.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__15384 (.I0(n10243), .I1(n10216), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5] ), 
            .I3(n10148), .O(n10244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__15384.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__15385 (.I0(n10229), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .O(n10245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__15385.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__15386 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[2] ), .O(n10246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15386.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15387 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[0] ), .O(n10247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f75 */ ;
    defparam LUT__15387.LUTMASK = 16'h1f75;
    EFX_LUT4 LUT__15388 (.I0(n10247), .I1(n10246), .I2(\i2c_config_index[4] ), 
            .I3(n10106), .O(n10248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__15388.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__15389 (.I0(n10248), .I1(n10245), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .O(n10249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15389.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15390 (.I0(n10243), .I1(n10171), .I2(n10230), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .O(n10250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8afc */ ;
    defparam LUT__15390.LUTMASK = 16'h8afc;
    EFX_LUT4 LUT__15391 (.I0(n10250), .I1(n10249), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__15391.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__15392 (.I0(n10251), .I1(n10244), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__15392.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__15393 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .O(n10252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15393.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15394 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .I2(n10151), .O(n10253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__15394.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__15395 (.I0(n10252), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6] ), 
            .I2(n10253), .I3(n10216), .O(n10254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__15395.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__15396 (.I0(\i2c_config_index[3] ), .I1(n10232), .I2(n10107), 
            .O(n10255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__15396.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__15397 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6] ), .I2(n10255), 
            .I3(n10161), .O(n10256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__15397.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__15398 (.I0(n10221), .I1(n10253), .I2(n10256), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077 */ ;
    defparam LUT__15398.LUTMASK = 16'hf077;
    EFX_LUT4 LUT__15399 (.I0(n10257), .I1(n10254), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15399.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15400 (.I0(n10243), .I1(n10151), .I2(\i2c_config_index[1] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), .O(n10258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ff5 */ ;
    defparam LUT__15400.LUTMASK = 16'h3ff5;
    EFX_LUT4 LUT__15401 (.I0(\i2c_config_index[2] ), .I1(n10258), .I2(n10142), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .O(n10259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15401.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15402 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7] ), .O(n10260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15402.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15403 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[3] ), .O(n10261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9ef3 */ ;
    defparam LUT__15403.LUTMASK = 16'h9ef3;
    EFX_LUT4 LUT__15404 (.I0(n10261), .I1(n10211), .I2(\i2c_config_index[4] ), 
            .I3(n10106), .O(n10262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__15404.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__15405 (.I0(n10262), .I1(n10260), .I2(n10161), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n10263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__15405.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__15406 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .I2(n10243), .O(n10264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__15406.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__15407 (.I0(n10252), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7] ), 
            .I2(n10264), .I3(n10216), .O(n10265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__15407.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__15408 (.I0(n10263), .I1(n10259), .I2(n10265), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__15408.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__15409 (.I0(\lcd_data[0] ), .I1(\lcd_data[1] ), .I2(\lcd_data[2] ), 
            .I3(\lcd_data[3] ), .O(n10266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6996 */ ;
    defparam LUT__15409.LUTMASK = 16'h6996;
    EFX_LUT4 LUT__15410 (.I0(\lcd_data[4] ), .I1(\lcd_data[3] ), .I2(n10266), 
            .O(n10267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15410.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15411 (.I0(\lcd_data[0] ), .I1(\lcd_data[1] ), .I2(\lcd_data[2] ), 
            .I3(\u_lcd_driver/n133 ), .O(n10268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he800 */ ;
    defparam LUT__15411.LUTMASK = 16'he800;
    EFX_LUT4 LUT__15412 (.I0(\u_lcd_driver/n133 ), .I1(\lcd_data[7] ), .O(n10269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15412.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15413 (.I0(\u_lcd_driver/n133 ), .I1(\lcd_data[5] ), .O(n10270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15413.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15414 (.I0(\lcd_data[3] ), .I1(\lcd_data[4] ), .I2(\u_lcd_driver/n133 ), 
            .O(n10271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__15414.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__15415 (.I0(\lcd_data[0] ), .I1(\lcd_data[1] ), .I2(\lcd_data[2] ), 
            .I3(\u_lcd_driver/n133 ), .O(n10272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9600 */ ;
    defparam LUT__15415.LUTMASK = 16'h9600;
    EFX_LUT4 LUT__15416 (.I0(\lcd_data[6] ), .I1(n10270), .I2(n10271), 
            .I3(n10272), .O(n10273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8ee8 */ ;
    defparam LUT__15416.LUTMASK = 16'h8ee8;
    EFX_LUT4 LUT__15417 (.I0(n10268), .I1(n10269), .I2(n10267), .I3(n10273), 
            .O(n10274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__15417.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__15418 (.I0(\lcd_data[5] ), .I1(\lcd_data[6] ), .I2(\u_lcd_driver/n133 ), 
            .O(n10275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__15418.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__15419 (.I0(n10272), .I1(n10271), .I2(n10275), .I3(n10269), 
            .O(n10276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9600 */ ;
    defparam LUT__15419.LUTMASK = 16'h9600;
    EFX_LUT4 LUT__15420 (.I0(\lcd_data[1] ), .I1(\lcd_data[3] ), .O(n10277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15420.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15421 (.I0(\lcd_data[2] ), .I1(\lcd_data[5] ), .I2(\lcd_data[6] ), 
            .I3(\lcd_data[7] ), .O(n10278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6996 */ ;
    defparam LUT__15421.LUTMASK = 16'h6996;
    EFX_LUT4 LUT__15422 (.I0(\lcd_data[0] ), .I1(\u_lcd_driver/n133 ), .O(n10279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15422.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15423 (.I0(\lcd_data[4] ), .I1(n10277), .I2(n10278), 
            .I3(n10279), .O(n10280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9600 */ ;
    defparam LUT__15423.LUTMASK = 16'h9600;
    EFX_LUT4 LUT__15424 (.I0(n10268), .I1(n10276), .I2(n10267), .I3(n10280), 
            .O(n10281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he8fe */ ;
    defparam LUT__15424.LUTMASK = 16'he8fe;
    EFX_LUT4 LUT__15425 (.I0(n10268), .I1(n10267), .I2(n10276), .I3(n10280), 
            .O(n10282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00e8 */ ;
    defparam LUT__15425.LUTMASK = 16'h00e8;
    EFX_LUT4 LUT__15426 (.I0(n10281), .I1(n10274), .I2(n10282), .O(n8110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__15426.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__15427 (.I0(n373), .I1(n366), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .O(n10283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15427.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15428 (.I0(n10272), .I1(n10271), .O(n10284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15428.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15429 (.I0(\lcd_data[4] ), .I1(n10277), .I2(n10266), 
            .I3(\u_lcd_driver/n133 ), .O(n10285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6000 */ ;
    defparam LUT__15429.LUTMASK = 16'h6000;
    EFX_LUT4 LUT__15430 (.I0(\lcd_data[0] ), .I1(\lcd_data[2] ), .O(n10286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15430.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15431 (.I0(n10274), .I1(n10281), .I2(n10282), .I3(n10286), 
            .O(n10287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bf4 */ ;
    defparam LUT__15431.LUTMASK = 16'h0bf4;
    EFX_LUT4 LUT__15432 (.I0(\lcd_data[4] ), .I1(n10277), .I2(n10286), 
            .O(n10288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7c7c */ ;
    defparam LUT__15432.LUTMASK = 16'h7c7c;
    EFX_LUT4 LUT__15433 (.I0(n10274), .I1(n10281), .I2(n10282), .I3(n10288), 
            .O(n10289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__15433.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__15434 (.I0(n10284), .I1(n10285), .I2(n10287), .I3(n10289), 
            .O(n10290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0017 */ ;
    defparam LUT__15434.LUTMASK = 16'h0017;
    EFX_LUT4 LUT__15435 (.I0(n10274), .I1(n10281), .I2(n10282), .I3(n10270), 
            .O(n10291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bf4 */ ;
    defparam LUT__15435.LUTMASK = 16'h0bf4;
    EFX_LUT4 LUT__15436 (.I0(n10277), .I1(n10291), .I2(n10275), .I3(n10284), 
            .O(n10292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h17e8 */ ;
    defparam LUT__15436.LUTMASK = 16'h17e8;
    EFX_LUT4 LUT__15437 (.I0(\lcd_data[0] ), .I1(\lcd_data[1] ), .I2(\u_lcd_driver/n133 ), 
            .O(n10293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__15437.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__15438 (.I0(n10272), .I1(n10279), .I2(n8110), .I3(n10293), 
            .O(n10294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he88e */ ;
    defparam LUT__15438.LUTMASK = 16'he88e;
    EFX_LUT4 LUT__15439 (.I0(\lcd_data[5] ), .I1(\lcd_data[7] ), .I2(n10277), 
            .I3(\u_lcd_driver/n133 ), .O(n8411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9600 */ ;
    defparam LUT__15439.LUTMASK = 16'h9600;
    EFX_LUT4 LUT__15440 (.I0(n10284), .I1(n10275), .O(n10295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15440.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15441 (.I0(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q ), .I1(\u_lcd_driver/r_lcd_dv~FF_frt_7_q ), 
            .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27_q ), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .O(n10296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4114 */ ;
    defparam LUT__15441.LUTMASK = 16'h4114;
    EFX_LUT4 LUT__15442 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q ), 
            .I1(n10296), .I2(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36_q ), 
            .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35_q ), .O(n10297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eef */ ;
    defparam LUT__15442.LUTMASK = 16'h8eef;
    EFX_LUT4 LUT__15443 (.I0(\u_rgb2dvi/enc_2/acc[0] ), .I1(\u_rgb2dvi/enc_2/acc[1] ), 
            .I2(\u_rgb2dvi/enc_2/acc[2] ), .I3(\u_rgb2dvi/enc_2/acc[3] ), 
            .O(n10298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15443.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15444 (.I0(\u_rgb2dvi/enc_2/acc[4] ), .I1(n10298), .O(n10299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15444.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15445 (.I0(n10297), .I1(n10299), .O(n10300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15445.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15446 (.I0(n387), .I1(n361), .I2(n10300), .O(n10301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15446.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15447 (.I0(n8411), .I1(n10269), .I2(n10295), .I3(n8110), 
            .O(n10302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1441 */ ;
    defparam LUT__15447.LUTMASK = 16'h1441;
    EFX_LUT4 LUT__15448 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38_q ), .I2(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36_q ), 
            .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35_q ), .O(n10303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd66b */ ;
    defparam LUT__15448.LUTMASK = 16'hd66b;
    EFX_LUT4 LUT__15449 (.I0(n10303), .I1(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q ), 
            .I2(\u_rgb2dvi/enc_2/acc[4] ), .I3(n10298), .O(n10304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__15449.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__15450 (.I0(n10301), .I1(n10283), .I2(n10304), .O(n5371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15450.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15451 (.I0(n362), .I1(n352), .I2(n10300), .O(n10305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15451.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15452 (.I0(n374), .I1(n367), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .O(n10306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15452.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15453 (.I0(n10306), .I1(n10305), .I2(n10304), .O(n5374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15453.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15454 (.I0(n388), .I1(n364), .I2(n10300), .O(n10307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15454.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15455 (.I0(n376), .I1(n369), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .O(n10308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15455.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15456 (.I0(n10308), .I1(n10307), .I2(n10304), .O(n5377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15456.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15457 (.I0(n3217), .I1(n3047), .I2(n10300), .O(n10309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15457.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15458 (.I0(n378), .I1(n371), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .O(n10310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15458.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15459 (.I0(n10310), .I1(n10309), .I2(n10304), .O(n5380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15459.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15460 (.I0(\u_rgb2dvi/enc_1/acc[0] ), .I1(\u_rgb2dvi/enc_1/acc[1] ), 
            .I2(\u_rgb2dvi/enc_1/acc[2] ), .I3(\u_rgb2dvi/enc_1/acc[3] ), 
            .O(n10311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15460.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15461 (.I0(\u_rgb2dvi/enc_1/acc[4] ), .I1(n10311), .O(n10312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15461.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15462 (.I0(n10297), .I1(n10312), .O(n10313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15462.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15463 (.I0(n387), .I1(n361), .I2(n10313), .O(n10314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15463.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15464 (.I0(n10303), .I1(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q ), 
            .I2(\u_rgb2dvi/enc_1/acc[4] ), .I3(n10311), .O(n10315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0ee */ ;
    defparam LUT__15464.LUTMASK = 16'he0ee;
    EFX_LUT4 LUT__15465 (.I0(n10314), .I1(n10283), .I2(n10315), .O(n5385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15465.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15466 (.I0(n362), .I1(n352), .I2(n10313), .O(n10316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15466.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15467 (.I0(n10316), .I1(n10306), .I2(n10315), .O(n5388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15467.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15468 (.I0(n388), .I1(n364), .I2(n10313), .O(n10317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15468.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15469 (.I0(n10317), .I1(n10308), .I2(n10315), .O(n5391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15469.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15470 (.I0(n3217), .I1(n3047), .I2(n10313), .O(n10318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15470.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15471 (.I0(n10318), .I1(n10310), .I2(n10315), .O(n5394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15471.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15472 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36_q ), .I2(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38_q ), 
            .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35_q ), .O(n5410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6996 */ ;
    defparam LUT__15472.LUTMASK = 16'h6996;
    EFX_LUT4 LUT__15473 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36_q ), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35_q ), 
            .I3(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38_q ), .O(n5416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdd4 */ ;
    defparam LUT__15473.LUTMASK = 16'hbdd4;
    EFX_LUT4 LUT__15474 (.I0(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q ), .I1(n5410), 
            .I2(n5416), .O(n5417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__15474.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__15475 (.I0(\u_lcd_driver/r_lcd_dv~FF_frt_7_q ), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27_q ), 
            .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), .O(n10319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__15475.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__15476 (.I0(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q ), .I1(n10319), 
            .I2(n5417), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q ), 
            .O(n5403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15476.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15477 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_37_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_6_frt_36_q ), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_35_q ), 
            .I3(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38_q ), .O(n5413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15477.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15478 (.I0(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q ), .I1(n5410), 
            .O(n5420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15478.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15479 (.I0(\u_rgb2dvi/enc_0/acc[4] ), .I1(n10297), .O(n10320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15479.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15480 (.I0(n387), .I1(n361), .I2(n10320), .O(n10321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15480.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15481 (.I0(\u_rgb2dvi/enc_0/acc[0] ), .I1(\u_rgb2dvi/enc_0/acc[1] ), 
            .I2(\u_rgb2dvi/enc_0/acc[2] ), .I3(\u_rgb2dvi/enc_0/acc[3] ), 
            .O(n10322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15481.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15482 (.I0(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q ), .I1(n10303), 
            .O(n10323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15482.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15483 (.I0(n10322), .I1(\u_rgb2dvi/enc_0/acc[4] ), .I2(n10323), 
            .O(n10324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__15483.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__15484 (.I0(n10321), .I1(n10283), .I2(n10324), .O(n5422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15484.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15485 (.I0(n362), .I1(n352), .I2(n10320), .O(n10325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15485.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15486 (.I0(n10325), .I1(n10306), .I2(n10324), .O(n5425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15486.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15487 (.I0(n388), .I1(n364), .I2(n10320), .O(n10326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15487.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15488 (.I0(n10326), .I1(n10308), .I2(n10324), .O(n5428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15488.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15489 (.I0(n3217), .I1(n3047), .I2(n10320), .O(n10327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15489.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15490 (.I0(n10327), .I1(n10310), .I2(n10324), .O(n5431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15490.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15493 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[0] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), 
            .O(\u_CMOS_Capture_RAW_Gray/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15493.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15494 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_href_r[1] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_href_r[0] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .O(ceg_net126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__15494.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__15496 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] ), 
            .O(\u_CMOS_Capture_RAW_Gray/n160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__15496.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__15497 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1] ), 
            .O(n10330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15497.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15498 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] ), 
            .I2(n10330), .O(ceg_net154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__15498.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__15499 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] ), 
            .I2(n10330), .O(\u_CMOS_Capture_RAW_Gray/n171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15499.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15530 (.I0(n445), .I1(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), 
            .O(\u_CMOS_Capture_RAW_Gray/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15530.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15531 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3236), 
            .O(\u_CMOS_Capture_RAW_Gray/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15531.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15532 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3234), 
            .O(\u_CMOS_Capture_RAW_Gray/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15532.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15533 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3232), 
            .O(\u_CMOS_Capture_RAW_Gray/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15533.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15534 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3230), 
            .O(\u_CMOS_Capture_RAW_Gray/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15534.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15535 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3228), 
            .O(\u_CMOS_Capture_RAW_Gray/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15535.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15536 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3226), 
            .O(\u_CMOS_Capture_RAW_Gray/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15536.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15537 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3224), 
            .O(\u_CMOS_Capture_RAW_Gray/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15537.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15538 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3222), 
            .O(\u_CMOS_Capture_RAW_Gray/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15538.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15539 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3220), 
            .O(\u_CMOS_Capture_RAW_Gray/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15539.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15540 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3219), 
            .O(\u_CMOS_Capture_RAW_Gray/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15540.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15541 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] ), 
            .O(\u_CMOS_Capture_RAW_Gray/n159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__15541.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__15577 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n5623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15577.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15578 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n5626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15578.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15579 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[1] ), .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[0] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/line_cnt[2] ), .I3(\u_CMOS_Capture_RAW_Gray/line_cnt[3] ), 
            .O(n10347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__15579.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__15580 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[4] ), .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[9] ), 
            .I2(n10347), .I3(\u_CMOS_Capture_RAW_Gray/line_cnt[8] ), .O(n10348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__15580.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__15581 (.I0(n10348), .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[5] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/line_cnt[8] ), .I3(\u_CMOS_Capture_RAW_Gray/line_cnt[9] ), 
            .O(n10349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf20d */ ;
    defparam LUT__15581.LUTMASK = 16'hf20d;
    EFX_LUT4 LUT__15582 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[8] ), .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[7] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/line_cnt[6] ), .I3(\u_CMOS_Capture_RAW_Gray/line_cnt[9] ), 
            .O(n10350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4001 */ ;
    defparam LUT__15582.LUTMASK = 16'h4001;
    EFX_LUT4 LUT__15583 (.I0(\u_CMOS_Capture_RAW_Gray/frame_sync_flag ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1] ), 
            .O(n10351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15583.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15584 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[10] ), .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[11] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/cmos_href_r[1] ), .I3(n10351), 
            .O(n10352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15584.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15585 (.I0(n10350), .I1(n10349), .I2(\u_CMOS_Capture_RAW_Gray/line_cnt[8] ), 
            .I3(n10352), .O(cmos_frame_href)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d00 */ ;
    defparam LUT__15585.LUTMASK = 16'h3d00;
    EFX_LUT4 LUT__15611 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n5660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15611.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15612 (.I0(\u_sensor_frame_count/delay_cnt[24] ), .I1(\u_sensor_frame_count/delay_cnt[25] ), 
            .O(n10353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15612.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15613 (.I0(\u_sensor_frame_count/delay_cnt[12] ), .I1(\u_sensor_frame_count/delay_cnt[26] ), 
            .I2(\u_sensor_frame_count/delay_cnt[16] ), .I3(\u_sensor_frame_count/delay_cnt[15] ), 
            .O(n10354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15613.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15614 (.I0(\u_sensor_frame_count/delay_cnt[0] ), .I1(\u_sensor_frame_count/delay_cnt[1] ), 
            .I2(\u_sensor_frame_count/delay_cnt[2] ), .I3(\u_sensor_frame_count/delay_cnt[5] ), 
            .O(n10355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15614.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15615 (.I0(\u_sensor_frame_count/delay_cnt[3] ), .I1(\u_sensor_frame_count/delay_cnt[4] ), 
            .I2(\u_sensor_frame_count/delay_cnt[6] ), .I3(\u_sensor_frame_count/delay_cnt[11] ), 
            .O(n10356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15615.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15616 (.I0(\u_sensor_frame_count/delay_cnt[7] ), .I1(\u_sensor_frame_count/delay_cnt[8] ), 
            .I2(\u_sensor_frame_count/delay_cnt[9] ), .I3(\u_sensor_frame_count/delay_cnt[10] ), 
            .O(n10357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15616.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15617 (.I0(n10355), .I1(n10356), .I2(n10357), .O(n10358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15617.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15618 (.I0(\u_sensor_frame_count/delay_cnt[14] ), .I1(\u_sensor_frame_count/delay_cnt[23] ), 
            .I2(\u_sensor_frame_count/delay_cnt[13] ), .I3(\u_sensor_frame_count/delay_cnt[27] ), 
            .O(n10359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15618.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15619 (.I0(\u_sensor_frame_count/delay_cnt[17] ), .I1(\u_sensor_frame_count/delay_cnt[18] ), 
            .I2(\u_sensor_frame_count/delay_cnt[19] ), .O(n10360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15619.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15620 (.I0(\u_sensor_frame_count/delay_cnt[20] ), .I1(\u_sensor_frame_count/delay_cnt[21] ), 
            .I2(\u_sensor_frame_count/delay_cnt[22] ), .O(n10361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15620.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15621 (.I0(n10359), .I1(n10360), .I2(n10361), .O(n10362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15621.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15622 (.I0(n10353), .I1(n10354), .I2(n10358), .I3(n10362), 
            .O(\u_sensor_frame_count/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__15622.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__15623 (.I0(\u_sensor_frame_count/cmos_fps_cnt[0] ), .I1(\u_sensor_frame_count/n110 ), 
            .O(\u_sensor_frame_count/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15623.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15624 (.I0(\u_sensor_frame_count/cmos_vsync_r[1] ), .I1(\u_sensor_frame_count/cmos_vsync_r[0] ), 
            .I2(\u_sensor_frame_count/n110 ), .O(ceg_net200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__15624.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__15625 (.I0(\u_scaler_gray/srcy_int[0] ), .I1(\u_scaler_gray/srcy_int[1] ), 
            .I2(\u_scaler_gray/srcy_int[2] ), .I3(\u_scaler_gray/srcy_int[3] ), 
            .O(n10363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15625.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15626 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] ), 
            .I1(\u_scaler_gray/srcy_int[5] ), .O(n10364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15626.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15627 (.I0(n10364), .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] ), 
            .I2(\u_scaler_gray/srcy_int[4] ), .I3(n10363), .O(n10365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7eeb */ ;
    defparam LUT__15627.LUTMASK = 16'h7eeb;
    EFX_LUT4 LUT__15628 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] ), 
            .I1(\u_scaler_gray/srcy_int[6] ), .O(n10366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15628.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15629 (.I0(\u_scaler_gray/srcy_int[4] ), .I1(\u_scaler_gray/srcy_int[5] ), 
            .I2(n10363), .O(n10367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15629.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15630 (.I0(n10366), .I1(n10367), .I2(n10365), .O(n10368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__15630.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__15631 (.I0(\u_scaler_gray/srcy_int[4] ), .I1(n10363), 
            .O(n10369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15631.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15632 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] ), 
            .I1(n10366), .I2(\u_scaler_gray/srcy_int[5] ), .I3(n10369), 
            .O(n10370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde */ ;
    defparam LUT__15632.LUTMASK = 16'hbdde;
    EFX_LUT4 LUT__15633 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] ), .I2(n10368), 
            .I3(n10370), .O(n10371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__15633.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__15634 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] ), 
            .I1(\u_scaler_gray/srcy_int[1] ), .I2(\u_scaler_gray/srcy_int[2] ), 
            .O(n10372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4 */ ;
    defparam LUT__15634.LUTMASK = 16'hd4d4;
    EFX_LUT4 LUT__15635 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] ), .I2(n10372), 
            .I3(\u_scaler_gray/srcy_int[3] ), .O(n10373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8ccf */ ;
    defparam LUT__15635.LUTMASK = 16'h8ccf;
    EFX_LUT4 LUT__15636 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] ), .I2(\u_scaler_gray/srcy_int[0] ), 
            .I3(\u_scaler_gray/srcy_int[1] ), .O(n10374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f75 */ ;
    defparam LUT__15636.LUTMASK = 16'h1f75;
    EFX_LUT4 LUT__15637 (.I0(\u_scaler_gray/srcy_int[0] ), .I1(\u_scaler_gray/srcy_int[1] ), 
            .O(n10375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15637.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15638 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] ), 
            .I1(\u_scaler_gray/srcy_int[3] ), .O(n10376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15638.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15639 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] ), 
            .I1(n10376), .I2(\u_scaler_gray/srcy_int[2] ), .I3(n10375), 
            .O(n10377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde */ ;
    defparam LUT__15639.LUTMASK = 16'hbdde;
    EFX_LUT4 LUT__15640 (.I0(n10377), .I1(n10374), .I2(n10363), .I3(n10373), 
            .O(n10378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__15640.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__15641 (.I0(n10378), .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] ), 
            .I2(n10370), .I3(n10368), .O(n10379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__15641.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__15642 (.I0(\u_scaler_gray/srcy_int[6] ), .I1(n10367), 
            .O(n10380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15642.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15643 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] ), 
            .I1(\u_scaler_gray/srcy_int[7] ), .I2(n10380), .O(n10381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__15643.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__15644 (.I0(\u_scaler_gray/srcy_int[4] ), .I1(\u_scaler_gray/srcy_int[5] ), 
            .O(n10382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15644.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15645 (.I0(\u_scaler_gray/srcy_int[6] ), .I1(\u_scaler_gray/srcy_int[7] ), 
            .I2(n10363), .I3(n10382), .O(n10383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15645.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15646 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] ), 
            .I1(\u_scaler_gray/srcy_int[9] ), .O(n10384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15646.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15647 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] ), 
            .I1(n10384), .I2(\u_scaler_gray/srcy_int[8] ), .I3(n10383), 
            .O(n10385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde */ ;
    defparam LUT__15647.LUTMASK = 16'hbdde;
    EFX_LUT4 LUT__15648 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] ), 
            .I1(\u_scaler_gray/srcy_int[7] ), .I2(n10380), .I3(n10385), 
            .O(n10386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__15648.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__15649 (.I0(n10379), .I1(n10381), .I2(n10371), .I3(n10386), 
            .O(n10387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__15649.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__15650 (.I0(\u_scaler_gray/srcy_int[8] ), .I1(\u_scaler_gray/srcy_int[9] ), 
            .O(n10388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15650.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15651 (.I0(\u_scaler_gray/srcy_int[6] ), .I1(\u_scaler_gray/srcy_int[7] ), 
            .I2(n10367), .I3(n10388), .O(n10389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15651.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15652 (.I0(\u_scaler_gray/srcy_int[10] ), .I1(n10389), 
            .O(n10390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__15652.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__15653 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] ), 
            .I1(\u_scaler_gray/srcy_int[8] ), .I2(n10383), .O(n10391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__15653.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__15654 (.I0(\u_scaler_gray/srcy_int[6] ), .I1(\u_scaler_gray/srcy_int[7] ), 
            .I2(\u_scaler_gray/srcy_int[8] ), .I3(n10367), .O(n10392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15654.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15655 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] ), 
            .I1(n10391), .I2(n10392), .I3(\u_scaler_gray/srcy_int[9] ), 
            .O(n10393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4dd4 */ ;
    defparam LUT__15655.LUTMASK = 16'h4dd4;
    EFX_LUT4 LUT__15656 (.I0(n10390), .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] ), 
            .I2(n10393), .O(n10394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__15656.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__15657 (.I0(\u_scaler_gray/srcy_int[10] ), .I1(n10389), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] ), .I3(\u_scaler_gray/srcy_int[11] ), 
            .O(n10395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8778 */ ;
    defparam LUT__15657.LUTMASK = 16'h8778;
    EFX_LUT4 LUT__15658 (.I0(\u_scaler_gray/srcy_int[10] ), .I1(\u_scaler_gray/srcy_int[11] ), 
            .I2(n10388), .O(n10396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15658.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15659 (.I0(n10383), .I1(n10396), .O(n10397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15659.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15660 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] ), 
            .I1(\u_scaler_gray/srcy_int[12] ), .I2(n10397), .O(n10398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__15660.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__15661 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] ), 
            .I1(n10390), .I2(n10395), .I3(n10398), .O(n10399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__15661.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__15662 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] ), 
            .I1(\u_scaler_gray/srcy_int[13] ), .O(n10400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15662.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15663 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] ), 
            .I1(\u_scaler_gray/srcy_int[12] ), .I2(n10397), .I3(n10400), 
            .O(n10401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3fd4 */ ;
    defparam LUT__15663.LUTMASK = 16'h3fd4;
    EFX_LUT4 LUT__15664 (.I0(n10398), .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] ), 
            .I2(n10395), .I3(n10401), .O(n10402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__15664.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__15665 (.I0(n10387), .I1(n10394), .I2(n10399), .I3(n10402), 
            .O(n10403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__15665.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__15666 (.I0(\u_scaler_gray/srcy_int[12] ), .I1(\u_scaler_gray/srcy_int[13] ), 
            .I2(n10383), .I3(n10396), .O(n10404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15666.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15667 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] ), 
            .I1(\u_scaler_gray/srcy_int[15] ), .O(n10405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15667.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15668 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] ), 
            .I1(n10405), .I2(\u_scaler_gray/srcy_int[14] ), .I3(n10404), 
            .O(n10406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde */ ;
    defparam LUT__15668.LUTMASK = 16'hbdde;
    EFX_LUT4 LUT__15669 (.I0(\u_scaler_gray/srcy_int[12] ), .I1(n10397), 
            .O(n10407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15669.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15670 (.I0(\u_scaler_gray/srcy_int[13] ), .I1(n10407), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] ), .O(n10408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__15670.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__15671 (.I0(n10406), .I1(n10408), .O(n10409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15671.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15672 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] ), 
            .I1(\u_scaler_gray/srcy_int[14] ), .I2(n10404), .O(n10410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4 */ ;
    defparam LUT__15672.LUTMASK = 16'hd4d4;
    EFX_LUT4 LUT__15673 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] ), 
            .I1(\u_scaler_gray/srcy_int[15] ), .I2(n10410), .O(n10411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4 */ ;
    defparam LUT__15673.LUTMASK = 16'hd4d4;
    EFX_LUT4 LUT__15674 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] ), .O(n10412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15674.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15675 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] ), .O(n10413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15675.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15676 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] ), .O(n10414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15676.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15677 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] ), .O(n10415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15677.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15678 (.I0(n10412), .I1(n10413), .I2(n10414), .I3(n10415), 
            .O(n10416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15678.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15679 (.I0(empty), .I1(n10416), .O(n10417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15679.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15680 (.I0(n10403), .I1(n10409), .I2(n10411), .I3(n10417), 
            .O(n197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__15680.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__15681 (.I0(n724), .I1(n2738), .I2(n2739), .I3(n2741), 
            .O(n10418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15681.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15682 (.I0(n2743), .I1(n2745), .I2(n2747), .I3(n2749), 
            .O(n10419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15682.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15683 (.I0(n2751), .I1(n2753), .I2(n2755), .I3(n2757), 
            .O(n10420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15683.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15684 (.I0(n2759), .I1(n2761), .I2(n2763), .O(n10421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15684.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15685 (.I0(n10418), .I1(n10419), .I2(n10420), .I3(n10421), 
            .O(n10422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15685.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15686 (.I0(n197), .I1(empty), .I2(n10422), .O(\u_afifo_buf/u_efx_fifo_top/rd_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__15686.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__15687 (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), .I1(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
            .O(n2090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15687.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15688 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[0] ), .I1(cmos_frame_href), 
            .O(\cmos_frame_Gray[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15688.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15689 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12] ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13] ), 
            .O(n10423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6996 */ ;
    defparam LUT__15689.LUTMASK = 16'h6996;
    EFX_LUT4 LUT__15690 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] ), 
            .I2(n10423), .O(n10424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__15690.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__15691 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3_q ), 
            .O(n10425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__15691.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__15692 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .I2(n10425), .O(n10426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__15692.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__15693 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .I2(n10426), .O(n10427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__15693.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__15694 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[2] ), .I1(n10427), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/waddr[1] ), .O(n10428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800 */ ;
    defparam LUT__15694.LUTMASK = 16'h1800;
    EFX_LUT4 LUT__15695 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[1] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[2] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] ), 
            .I3(n10427), .O(n10429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4001 */ ;
    defparam LUT__15695.LUTMASK = 16'h4001;
    EFX_LUT4 LUT__15696 (.I0(n10428), .I1(n10429), .I2(\u_afifo_buf/u_efx_fifo_top/waddr[0] ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] ), 
            .O(n10430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaac */ ;
    defparam LUT__15696.LUTMASK = 16'hcaac;
    EFX_LUT4 LUT__15697 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[5] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[6] ), 
            .I2(n10425), .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .O(n10431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbd7e */ ;
    defparam LUT__15697.LUTMASK = 16'hbd7e;
    EFX_LUT4 LUT__15698 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[3] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[4] ), 
            .I2(n10426), .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .O(n10432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbd7e */ ;
    defparam LUT__15698.LUTMASK = 16'hbd7e;
    EFX_LUT4 LUT__15699 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[7] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[8] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF_frt_3_q ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .O(n10433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbd7e */ ;
    defparam LUT__15699.LUTMASK = 16'hbd7e;
    EFX_LUT4 LUT__15700 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[9] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[10] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2_q ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] ), 
            .O(n10434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbd7e */ ;
    defparam LUT__15700.LUTMASK = 16'hbd7e;
    EFX_LUT4 LUT__15701 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13] ), 
            .O(n10435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15701.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15702 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[11] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), 
            .I2(n10435), .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] ), 
            .O(n10436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbd7e */ ;
    defparam LUT__15702.LUTMASK = 16'hbd7e;
    EFX_LUT4 LUT__15703 (.I0(n10434), .I1(n10436), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13] ), 
            .O(n10437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110 */ ;
    defparam LUT__15703.LUTMASK = 16'h0110;
    EFX_LUT4 LUT__15704 (.I0(n10431), .I1(n10432), .I2(n10433), .I3(n10437), 
            .O(n10438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15704.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15705 (.I0(n10438), .I1(n10430), .I2(cmos_frame_href), 
            .O(\u_afifo_buf/u_efx_fifo_top/wr_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__15705.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__15706 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), .I1(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15706.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15707 (.I0(\u_sensor_frame_count/delay_cnt[12] ), .I1(n10358), 
            .I2(\u_sensor_frame_count/delay_cnt[13] ), .I3(\u_sensor_frame_count/delay_cnt[14] ), 
            .O(n10439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__15707.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__15708 (.I0(n10439), .I1(\u_sensor_frame_count/delay_cnt[15] ), 
            .I2(\u_sensor_frame_count/delay_cnt[16] ), .I3(n10360), .O(n10440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__15708.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__15709 (.I0(n10440), .I1(n10361), .I2(\u_sensor_frame_count/delay_cnt[23] ), 
            .I3(n10353), .O(n10441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__15709.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__15710 (.I0(n10441), .I1(\u_sensor_frame_count/delay_cnt[26] ), 
            .I2(\u_sensor_frame_count/delay_cnt[27] ), .O(n10442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__15710.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__15711 (.I0(\u_sensor_frame_count/delay_cnt[0] ), .I1(n10442), 
            .O(\u_sensor_frame_count/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15711.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15712 (.I0(n10442), .I1(n575), .O(\u_sensor_frame_count/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15712.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15713 (.I0(n10442), .I1(n3091), .O(\u_sensor_frame_count/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15713.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15714 (.I0(n10442), .I1(n3089), .O(\u_sensor_frame_count/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15714.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15715 (.I0(n10442), .I1(n3087), .O(\u_sensor_frame_count/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15715.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15716 (.I0(n10442), .I1(n3085), .O(\u_sensor_frame_count/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15716.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15717 (.I0(n10442), .I1(n3083), .O(\u_sensor_frame_count/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15717.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15718 (.I0(n10442), .I1(n3081), .O(\u_sensor_frame_count/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15718.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15719 (.I0(n10442), .I1(n3079), .O(\u_sensor_frame_count/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15719.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15720 (.I0(n10442), .I1(n3077), .O(\u_sensor_frame_count/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15720.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15721 (.I0(n10442), .I1(n3075), .O(\u_sensor_frame_count/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15721.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15722 (.I0(n10442), .I1(n3062), .O(\u_sensor_frame_count/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15722.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15723 (.I0(n10442), .I1(n3060), .O(\u_sensor_frame_count/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15723.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15724 (.I0(n10442), .I1(n3055), .O(\u_sensor_frame_count/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15724.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15725 (.I0(n10442), .I1(n3053), .O(\u_sensor_frame_count/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15725.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15726 (.I0(n10442), .I1(n3049), .O(\u_sensor_frame_count/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15726.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15727 (.I0(n10442), .I1(n3045), .O(\u_sensor_frame_count/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15727.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15728 (.I0(n10442), .I1(n3041), .O(\u_sensor_frame_count/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15728.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15729 (.I0(n10442), .I1(n2910), .O(\u_sensor_frame_count/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15729.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15730 (.I0(n10442), .I1(n2908), .O(\u_sensor_frame_count/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15730.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15731 (.I0(n10442), .I1(n2891), .O(\u_sensor_frame_count/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15731.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15732 (.I0(n10442), .I1(n2889), .O(\u_sensor_frame_count/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15732.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15733 (.I0(n10442), .I1(n2887), .O(\u_sensor_frame_count/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15733.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15734 (.I0(n10442), .I1(n2885), .O(\u_sensor_frame_count/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15734.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15735 (.I0(n10442), .I1(n2883), .O(\u_sensor_frame_count/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15735.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15736 (.I0(n10442), .I1(n2881), .O(\u_sensor_frame_count/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15736.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15737 (.I0(n10442), .I1(n2879), .O(\u_sensor_frame_count/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15737.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15738 (.I0(n10442), .I1(n2878), .O(\u_sensor_frame_count/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15738.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15739 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n5723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15739.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15740 (.I0(n601), .I1(\u_sensor_frame_count/n110 ), .O(\u_sensor_frame_count/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15740.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15741 (.I0(n2876), .I1(\u_sensor_frame_count/n110 ), .O(\u_sensor_frame_count/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15741.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15742 (.I0(n2874), .I1(\u_sensor_frame_count/n110 ), .O(\u_sensor_frame_count/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15742.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15743 (.I0(n2872), .I1(\u_sensor_frame_count/n110 ), .O(\u_sensor_frame_count/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15743.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15744 (.I0(n2870), .I1(\u_sensor_frame_count/n110 ), .O(\u_sensor_frame_count/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15744.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15745 (.I0(n2868), .I1(\u_sensor_frame_count/n110 ), .O(\u_sensor_frame_count/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15745.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15746 (.I0(n2866), .I1(\u_sensor_frame_count/n110 ), .O(\u_sensor_frame_count/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15746.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15747 (.I0(n2865), .I1(\u_sensor_frame_count/n110 ), .O(\u_sensor_frame_count/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15747.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15748 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n5734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15748.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15749 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n5737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15749.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15750 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n5740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__15750.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__15751 (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), .I1(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
            .O(n2104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15751.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15752 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[2] ), .I1(cmos_frame_href), 
            .O(\cmos_frame_Gray[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15752.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15753 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), .I1(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15753.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15754 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[1] ), .I1(cmos_frame_href), 
            .O(\cmos_frame_Gray[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15754.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15755 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[3] ), .I1(cmos_frame_href), 
            .O(\cmos_frame_Gray[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15755.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15756 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[4] ), .I1(cmos_frame_href), 
            .O(\cmos_frame_Gray[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15756.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15757 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[5] ), .I1(cmos_frame_href), 
            .O(\cmos_frame_Gray[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15757.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15758 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[6] ), .I1(cmos_frame_href), 
            .O(\cmos_frame_Gray[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15758.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15759 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[7] ), .I1(cmos_frame_href), 
            .O(\cmos_frame_Gray[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15759.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15760 (.I0(n10422), .I1(empty), .I2(n197), .O(ceg_net219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15760.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15761 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13] ), 
            .O(n7826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15761.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15762 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11] ), 
            .I1(n7826), .O(n7829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15762.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15763 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF_frt_1_q ), 
            .O(n7832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15763.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15764 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] ), 
            .I1(n7832), .O(n7835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15764.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15765 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .I1(n7835), .O(n7838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15765.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15766 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .I3(n7838), .O(n7847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6996 */ ;
    defparam LUT__15766.LUTMASK = 16'h6996;
    EFX_LUT4 LUT__15767 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .I1(n7847), .O(n7850)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15767.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15768 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .I2(n7850), .O(n7856)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__15768.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__15769 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] ), 
            .I2(n7856), .O(n5807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__15769.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__15770 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .O(n10443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15770.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15771 (.I0(n10443), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[0] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[1] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15771.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15772 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[0] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[1] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15772.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15775 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .O(n10444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15775.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15776 (.I0(n10444), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[1] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[2] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15776.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15777 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .O(n10445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15777.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15778 (.I0(n10445), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[2] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[3] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15778.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15779 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .O(n10446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15779.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15780 (.I0(n10446), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[3] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[4] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15780.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15781 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .O(n10447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15781.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15782 (.I0(n10447), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[4] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[5] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15782.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15783 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .O(n10448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15783.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15784 (.I0(n10448), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[5] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[6] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15784.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15785 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .O(n10449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15785.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15786 (.I0(n10449), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[6] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[7] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15786.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15787 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .O(n10450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15787.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15788 (.I0(n10450), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[7] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[8] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15788.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15789 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .O(n10451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15789.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15790 (.I0(n10451), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[8] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[9] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15790.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15791 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] ), 
            .O(n10452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15791.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15792 (.I0(n10452), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[9] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[10] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15792.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15793 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] ), 
            .O(n10453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15793.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15794 (.I0(n10453), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[10] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[11] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__15794.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__15795 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), .I2(empty), .O(n10454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15795.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15796 (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[11] ), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] ), 
            .I2(empty), .I3(n10454), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h53ac */ ;
    defparam LUT__15796.LUTMASK = 16'h53ac;
    EFX_LUT4 LUT__15797 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] ), 
            .I2(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15797.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15798 (.I0(n10454), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[13] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15798.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15799 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[1] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[2] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15799.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15800 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[2] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[3] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15800.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15801 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[3] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[4] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15801.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15802 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[4] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[5] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15802.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15803 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[5] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[6] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15803.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15804 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[6] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[7] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15804.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15805 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[7] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[8] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15805.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15806 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[8] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[9] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15806.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15807 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[9] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[10] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15807.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15808 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[10] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[11] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15808.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15809 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[11] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15809.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15810 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15810.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15811 (.I0(tvalid_o), .I1(\u_scaler_gray/tvalid_o_r ), 
            .O(ceg_net226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__15811.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__15812 (.I0(\u_scaler_gray/vs_cnt[12] ), .I1(\u_scaler_gray/vs_cnt[13] ), 
            .I2(\u_scaler_gray/vs_cnt[14] ), .I3(\u_scaler_gray/vs_cnt[15] ), 
            .O(n10455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15812.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15813 (.I0(\u_scaler_gray/vs_cnt[3] ), .I1(\u_scaler_gray/vs_cnt[5] ), 
            .I2(\u_scaler_gray/vs_cnt[7] ), .I3(\u_scaler_gray/vs_cnt[8] ), 
            .O(n10456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15813.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15814 (.I0(\u_scaler_gray/vs_cnt[10] ), .I1(\u_scaler_gray/vs_cnt[11] ), 
            .I2(n10455), .I3(n10456), .O(n10457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15814.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15815 (.I0(\u_scaler_gray/vs_cnt[0] ), .I1(\u_scaler_gray/vs_cnt[6] ), 
            .I2(\u_scaler_gray/vs_cnt[9] ), .I3(tvalid_o), .O(n10458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15815.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15816 (.I0(\u_scaler_gray/tvalid_o_r ), .I1(\u_scaler_gray/vs_cnt[1] ), 
            .I2(\u_scaler_gray/vs_cnt[2] ), .I3(\u_scaler_gray/vs_cnt[4] ), 
            .O(n10459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15816.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15817 (.I0(n10457), .I1(n10458), .I2(n10459), .O(\u_scaler_gray/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15817.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15818 (.I0(\u_scaler_gray/vs_cnt[2] ), .I1(\u_scaler_gray/vs_cnt[4] ), 
            .I2(\u_scaler_gray/vs_cnt[6] ), .I3(\u_scaler_gray/vs_cnt[9] ), 
            .O(n10460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15818.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15819 (.I0(ceg_net226), .I1(\u_scaler_gray/vs_cnt[1] ), 
            .I2(\u_scaler_gray/vs_cnt[0] ), .O(n10461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__15819.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__15820 (.I0(n10457), .I1(n10460), .I2(n10461), .O(n10462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15820.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15821 (.I0(\u_scaler_gray/n150 ), .I1(n10462), .O(ceg_net229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__15821.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__15822 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1] ), .O(n10463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15822.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15823 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7] ), .O(n10464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15823.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15824 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0] ), .O(n10465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15824.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15825 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15] ), .O(n10466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15825.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15826 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10] ), .I2(n10465), 
            .I3(n10466), .O(n10467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__15826.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__15827 (.I0(n197), .I1(n10463), .I2(n10464), .I3(n10467), 
            .O(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15827.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15828 (.I0(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .I3(\Axi0ResetReg[2] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1703 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h80ff */ ;
    defparam LUT__15828.LUTMASK = 16'h80ff;
    EFX_LUT4 LUT__15829 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[12] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_addra[13] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_addra[14] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_addra[15] ), .O(n10468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15829.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15830 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[9] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_addra[10] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_addra[0] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_addra[11] ), .O(n10469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15830.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15831 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[4] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_addra[5] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_addra[6] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_addra[7] ), .O(n10470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15831.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15832 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_addra[2] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_addra[3] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_addra[8] ), .O(n10471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15832.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15833 (.I0(n10468), .I1(n10469), .I2(n10470), .I3(n10471), 
            .O(n10472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15833.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15834 (.I0(n197), .I1(n10472), .I2(\Axi0ResetReg[2] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1704 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f */ ;
    defparam LUT__15834.LUTMASK = 16'h8f8f;
    EFX_LUT4 LUT__15835 (.I0(\u_scaler_gray/srcy_int[12] ), .I1(\u_scaler_gray/srcy_int[13] ), 
            .I2(\u_scaler_gray/srcy_int[14] ), .I3(\u_scaler_gray/srcy_int[15] ), 
            .O(n10473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15835.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15836 (.I0(\u_scaler_gray/srcy_int[8] ), .I1(\u_scaler_gray/srcy_int[10] ), 
            .I2(\u_scaler_gray/srcy_int[11] ), .I3(\u_scaler_gray/srcy_int[9] ), 
            .O(n10474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15836.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15837 (.I0(\u_scaler_gray/srcy_int[4] ), .I1(\u_scaler_gray/srcy_int[5] ), 
            .I2(\u_scaler_gray/srcy_int[6] ), .I3(\u_scaler_gray/srcy_int[7] ), 
            .O(n10475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15837.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15838 (.I0(n10363), .I1(n10473), .I2(n10474), .I3(n10475), 
            .O(n10476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15838.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15839 (.I0(n10403), .I1(n10409), .I2(n10411), .O(n10477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__15839.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__15840 (.I0(\u_scaler_gray/destx[10] ), .I1(\u_scaler_gray/destx[11] ), 
            .I2(\u_scaler_gray/destx[8] ), .I3(\u_scaler_gray/destx[9] ), 
            .O(n10478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15840.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15841 (.I0(\u_scaler_gray/destx[12] ), .I1(\u_scaler_gray/destx[13] ), 
            .I2(\u_scaler_gray/destx[14] ), .I3(\u_scaler_gray/destx[15] ), 
            .O(n10479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15841.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15842 (.I0(\u_scaler_gray/destx[0] ), .I1(\u_scaler_gray/destx[1] ), 
            .I2(\u_scaler_gray/destx[2] ), .I3(\u_scaler_gray/destx[3] ), 
            .O(n10480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15842.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15843 (.I0(\u_scaler_gray/destx[4] ), .I1(\u_scaler_gray/destx[5] ), 
            .I2(\u_scaler_gray/destx[6] ), .I3(\u_scaler_gray/destx[7] ), 
            .O(n10481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15843.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15844 (.I0(n10478), .I1(n10479), .I2(n10480), .I3(n10481), 
            .O(n10482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15844.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15845 (.I0(n10477), .I1(n10476), .I2(n10482), .I3(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), 
            .O(n10483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__15845.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__15846 (.I0(n10416), .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), .I3(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), 
            .O(n10484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc700 */ ;
    defparam LUT__15846.LUTMASK = 16'hc700;
    EFX_LUT4 LUT__15847 (.I0(\u_scaler_gray/desty[12] ), .I1(\u_scaler_gray/desty[13] ), 
            .I2(\u_scaler_gray/desty[14] ), .I3(\u_scaler_gray/desty[15] ), 
            .O(n10485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15847.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15848 (.I0(\u_scaler_gray/desty[3] ), .I1(\u_scaler_gray/desty[5] ), 
            .I2(\u_scaler_gray/desty[7] ), .I3(\u_scaler_gray/desty[8] ), 
            .O(n10486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15848.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15849 (.I0(\u_scaler_gray/desty[10] ), .I1(\u_scaler_gray/desty[11] ), 
            .I2(n10485), .I3(n10486), .O(n10487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15849.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15850 (.I0(\u_scaler_gray/desty[2] ), .I1(\u_scaler_gray/desty[4] ), 
            .I2(\u_scaler_gray/desty[6] ), .I3(\u_scaler_gray/desty[9] ), 
            .O(n10488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15850.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15851 (.I0(\u_scaler_gray/desty[0] ), .I1(\u_scaler_gray/desty[1] ), 
            .I2(n10487), .I3(n10488), .O(n10489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15851.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15852 (.I0(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[0] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[1] ), .I2(n10489), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), .O(n10490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__15852.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__15853 (.I0(n10490), .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), .O(n10491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__15853.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__15854 (.I0(n10483), .I1(n10484), .I2(n10491), .I3(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h03ac */ ;
    defparam LUT__15854.LUTMASK = 16'h03ac;
    EFX_LUT4 LUT__15855 (.I0(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[0] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), .O(\u_scaler_gray/u0_data_stream_ctr/n2157 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15855.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15856 (.I0(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .I3(\Axi0ResetReg[2] ), .O(ceg_net526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbeaa */ ;
    defparam LUT__15856.LUTMASK = 16'hbeaa;
    EFX_LUT4 LUT__15857 (.I0(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__15857.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__15858 (.I0(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
            .I1(n10482), .O(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15858.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15859 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
            .I1(\Axi0ResetReg[2] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__15859.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__15860 (.I0(\u_scaler_gray/desty[0] ), .I1(\u_scaler_gray/desty[1] ), 
            .I2(\u_scaler_gray/desty[2] ), .I3(\u_scaler_gray/desty[4] ), 
            .O(n10492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15860.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15861 (.I0(\u_scaler_gray/desty[6] ), .I1(\u_scaler_gray/desty[9] ), 
            .I2(n10487), .I3(n10492), .O(n10493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15861.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15862 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
            .I1(n10493), .I2(\Axi0ResetReg[2] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1713 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f */ ;
    defparam LUT__15862.LUTMASK = 16'h8f8f;
    EFX_LUT4 LUT__15863 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n87 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n86 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15863.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15864 (.I0(\u_scaler_gray/srcx_int[4] ), .I1(\u_scaler_gray/srcx_int[5] ), 
            .I2(\u_scaler_gray/srcx_int[6] ), .I3(\u_scaler_gray/srcx_int[7] ), 
            .O(n10494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15864.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15865 (.I0(\u_scaler_gray/srcx_int[0] ), .I1(\u_scaler_gray/srcx_int[1] ), 
            .I2(\u_scaler_gray/srcx_int[2] ), .I3(\u_scaler_gray/srcx_int[3] ), 
            .O(n10495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15865.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15866 (.I0(n10494), .I1(n10495), .O(n10496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15866.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15867 (.I0(\u_scaler_gray/srcx_int[12] ), .I1(\u_scaler_gray/srcx_int[13] ), 
            .I2(\u_scaler_gray/srcx_int[14] ), .I3(\u_scaler_gray/srcx_int[15] ), 
            .O(n10497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15867.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15868 (.I0(\u_scaler_gray/srcx_int[8] ), .I1(\u_scaler_gray/srcx_int[9] ), 
            .I2(\u_scaler_gray/srcx_int[11] ), .I3(\u_scaler_gray/srcx_int[10] ), 
            .O(n10498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__15868.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__15869 (.I0(n10497), .I1(n10498), .O(n10499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15869.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15870 (.I0(n10499), .I1(n10496), .I2(\u_scaler_gray/srcx_int[0] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n903 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__15870.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__15871 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n102 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n101 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15871.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15872 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), 
            .I1(\Axi0ResetReg[2] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1702 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__15872.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__15873 (.I0(n10491), .I1(n10484), .I2(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf1f1 */ ;
    defparam LUT__15873.LUTMASK = 16'hf1f1;
    EFX_LUT4 LUT__15874 (.I0(n10489), .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), .I3(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ecc */ ;
    defparam LUT__15874.LUTMASK = 16'h0ecc;
    EFX_LUT4 LUT__15875 (.I0(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[0] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[1] ), .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n2080 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__15875.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__15876 (.I0(\u_scaler_gray/srcx_int[8] ), .I1(\u_scaler_gray/srcy_int[0] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15876.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15877 (.I0(\u_scaler_gray/srcx_int[8] ), .I1(\u_scaler_gray/srcy_int[0] ), 
            .I2(\u_scaler_gray/srcx_int[9] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__15877.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__15878 (.I0(\u_scaler_gray/srcx_int[8] ), .I1(\u_scaler_gray/srcx_int[9] ), 
            .O(n10500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15878.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15879 (.I0(n10500), .I1(\u_scaler_gray/srcy_int[0] ), 
            .I2(\u_scaler_gray/srcx_int[10] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__15879.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__15880 (.I0(\u_scaler_gray/srcx_int[10] ), .I1(n10500), 
            .I2(\u_scaler_gray/srcy_int[0] ), .I3(\u_scaler_gray/srcx_int[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1fe0 */ ;
    defparam LUT__15880.LUTMASK = 16'h1fe0;
    EFX_LUT4 LUT__15881 (.I0(\u_scaler_gray/srcx_int[1] ), .I1(\u_scaler_gray/u0_data_stream_ctr/n903 ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n885 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15881.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15882 (.I0(\u_scaler_gray/srcx_int[1] ), .I1(\u_scaler_gray/u0_data_stream_ctr/n903 ), 
            .I2(\u_scaler_gray/srcx_int[2] ), .O(\u_scaler_gray/u0_data_stream_ctr/n884 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__15882.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__15883 (.I0(\u_scaler_gray/srcx_int[1] ), .I1(\u_scaler_gray/srcx_int[2] ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/n903 ), .I3(\u_scaler_gray/srcx_int[3] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n883 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__15883.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__15884 (.I0(n10499), .I1(n10496), .I2(n10495), .O(n10501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__15884.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__15885 (.I0(\u_scaler_gray/srcx_int[4] ), .I1(n10501), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n882 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15885.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15886 (.I0(\u_scaler_gray/srcx_int[4] ), .I1(n10501), 
            .O(n10502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15886.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15887 (.I0(\u_scaler_gray/srcx_int[5] ), .I1(n10502), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n881 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15887.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15888 (.I0(\u_scaler_gray/srcx_int[5] ), .I1(n10502), 
            .I2(\u_scaler_gray/srcx_int[6] ), .O(\u_scaler_gray/u0_data_stream_ctr/n880 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__15888.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__15889 (.I0(\u_scaler_gray/srcx_int[5] ), .I1(\u_scaler_gray/srcx_int[6] ), 
            .I2(n10502), .I3(\u_scaler_gray/srcx_int[7] ), .O(\u_scaler_gray/u0_data_stream_ctr/n879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__15889.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__15890 (.I0(n10499), .I1(n10496), .O(n10503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15890.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15891 (.I0(\u_scaler_gray/u0_data_stream_ctr/n1162 ), .I1(n10503), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15891.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15892 (.I0(\u_scaler_gray/srcx_int[8] ), .I1(\u_scaler_gray/srcy_int[0] ), 
            .I2(n10503), .I3(\u_scaler_gray/srcx_int[9] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h17e8 */ ;
    defparam LUT__15892.LUTMASK = 16'h17e8;
    EFX_LUT4 LUT__15893 (.I0(\u_scaler_gray/srcx_int[9] ), .I1(\u_scaler_gray/srcx_int[8] ), 
            .I2(n10496), .I3(\u_scaler_gray/srcy_int[0] ), .O(n10504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha87f */ ;
    defparam LUT__15893.LUTMASK = 16'ha87f;
    EFX_LUT4 LUT__15894 (.I0(\u_scaler_gray/srcx_int[10] ), .I1(n10504), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__15894.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__15895 (.I0(\u_scaler_gray/srcx_int[10] ), .I1(\u_scaler_gray/srcy_int[0] ), 
            .I2(\u_scaler_gray/srcx_int[11] ), .I3(n10504), .O(\u_scaler_gray/u0_data_stream_ctr/n1176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3c5a */ ;
    defparam LUT__15895.LUTMASK = 16'h3c5a;
    EFX_LUT4 LUT__15896 (.I0(\u_scaler_gray/srcy_int[0] ), .I1(\u_scaler_gray/srcx_int[8] ), 
            .I2(\u_scaler_gray/srcx_int[9] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1195 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__15896.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__15897 (.I0(\u_scaler_gray/srcy_int[0] ), .I1(n10500), 
            .I2(\u_scaler_gray/srcx_int[10] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1e1 */ ;
    defparam LUT__15897.LUTMASK = 16'he1e1;
    EFX_LUT4 LUT__15898 (.I0(\u_scaler_gray/srcx_int[10] ), .I1(n10500), 
            .I2(\u_scaler_gray/srcy_int[0] ), .I3(\u_scaler_gray/srcx_int[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf10e */ ;
    defparam LUT__15898.LUTMASK = 16'hf10e;
    EFX_LUT4 LUT__15899 (.I0(\u_scaler_gray/srcx_int[8] ), .I1(\u_scaler_gray/srcy_int[0] ), 
            .I2(n10503), .I3(\u_scaler_gray/srcx_int[9] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1212 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4db2 */ ;
    defparam LUT__15899.LUTMASK = 16'h4db2;
    EFX_LUT4 LUT__15900 (.I0(\u_scaler_gray/srcx_int[9] ), .I1(\u_scaler_gray/srcx_int[8] ), 
            .I2(n10496), .I3(\u_scaler_gray/srcy_int[0] ), .O(n10505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fa8 */ ;
    defparam LUT__15900.LUTMASK = 16'h7fa8;
    EFX_LUT4 LUT__15901 (.I0(\u_scaler_gray/srcx_int[10] ), .I1(n10505), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1211 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__15901.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__15902 (.I0(\u_scaler_gray/srcx_int[10] ), .I1(\u_scaler_gray/srcy_int[0] ), 
            .I2(\u_scaler_gray/srcx_int[11] ), .I3(n10505), .O(\u_scaler_gray/u0_data_stream_ctr/n1210 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc35a */ ;
    defparam LUT__15902.LUTMASK = 16'hc35a;
    EFX_LUT4 LUT__15903 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n90 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n89 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15903.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15904 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n84 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n83 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15904.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15905 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n93 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n92 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15905.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15906 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n99 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n98 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15906.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15907 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n96 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n95 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15907.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15908 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n104 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n105 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15908.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15909 (.I0(n10462), .I1(n745), .O(\u_scaler_gray/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15909.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15910 (.I0(n10462), .I1(n2702), .O(\u_scaler_gray/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15910.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15911 (.I0(n10462), .I1(n2700), .O(\u_scaler_gray/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15911.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15912 (.I0(n10462), .I1(n2696), .O(\u_scaler_gray/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15912.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15913 (.I0(n10462), .I1(n2694), .O(\u_scaler_gray/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15913.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15914 (.I0(n10462), .I1(n2691), .O(\u_scaler_gray/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15914.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15915 (.I0(n10462), .I1(n2689), .O(\u_scaler_gray/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15915.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15916 (.I0(n10462), .I1(n2687), .O(\u_scaler_gray/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15916.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15917 (.I0(n10462), .I1(n2605), .O(\u_scaler_gray/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15917.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15918 (.I0(n10462), .I1(n2603), .O(\u_scaler_gray/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15918.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15919 (.I0(n10462), .I1(n2601), .O(\u_scaler_gray/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15919.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15920 (.I0(n10462), .I1(n2599), .O(\u_scaler_gray/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15920.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15921 (.I0(n10462), .I1(n2597), .O(\u_scaler_gray/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15921.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15922 (.I0(n10462), .I1(n2595), .O(\u_scaler_gray/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15922.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15923 (.I0(n10462), .I1(n2594), .O(\u_scaler_gray/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__15923.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__15924 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15] ), 
            .O(n10506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15924.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15925 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26] ), 
            .O(n10507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15925.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15926 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27] ), 
            .O(n10508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15926.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15927 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23] ), 
            .O(n10509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15927.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15928 (.I0(n10507), .I1(n10508), .I2(n10509), .O(n10510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15928.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15929 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18] ), 
            .I2(n10506), .I3(n10510), .O(n10511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15929.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15930 (.I0(n1656), .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0] ), 
            .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15930.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15931 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15] ), 
            .O(n10512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15931.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15932 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26] ), 
            .O(n10513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__15932.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__15933 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27] ), 
            .O(n10514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15933.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15934 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23] ), 
            .O(n10515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__15934.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__15935 (.I0(n10513), .I1(n10514), .I2(n10515), .O(n10516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__15935.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__15936 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18] ), 
            .I2(n10512), .I3(n10516), .O(n10517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__15936.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__15937 (.I0(DdrCtrl_ALEN_0[0]), .I1(n1487), .I2(n10517), 
            .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15937.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15938 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10] ), 
            .I1(n1485), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15938.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15939 (.I0(n1654), .I1(n1483), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n333 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15939.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15940 (.I0(n1481), .I1(n1371), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15940.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15941 (.I0(n1479), .I1(n1369), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15941.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15942 (.I0(n1477), .I1(n1367), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15942.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15943 (.I0(n1475), .I1(n1365), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n329 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15943.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15944 (.I0(n1473), .I1(n1363), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15944.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15945 (.I0(n1471), .I1(n1339), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n327 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15945.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15946 (.I0(n1469), .I1(n1337), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15946.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15947 (.I0(n1467), .I1(n1335), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15947.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15948 (.I0(n1465), .I1(n1333), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15948.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15949 (.I0(n1463), .I1(n1331), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n323 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15949.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15950 (.I0(n1419), .I1(n1329), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15950.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15951 (.I0(n1417), .I1(n1327), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n321 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15951.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15952 (.I0(n1415), .I1(n1325), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15952.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15953 (.I0(n1413), .I1(n1323), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15953.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15954 (.I0(n1411), .I1(n1321), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15954.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15955 (.I0(n1410), .I1(n1320), .I2(n10517), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15955.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15956 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1] ), 
            .I1(n1318), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15956.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15957 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2] ), 
            .I1(n1316), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15957.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15958 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3] ), 
            .I1(n1314), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15958.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15959 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4] ), 
            .I1(n1312), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15959.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15960 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5] ), 
            .I1(n1310), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15960.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15961 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6] ), 
            .I1(n1308), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15961.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15962 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7] ), 
            .I1(n1306), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15962.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15963 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8] ), 
            .I1(n1304), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15963.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15964 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9] ), 
            .I1(n1302), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15964.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15965 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10] ), 
            .I1(n1300), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15965.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15966 (.I0(n1686), .I1(n1298), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15966.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15967 (.I0(n1296), .I1(n1261), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15967.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15968 (.I0(n1294), .I1(n1259), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15968.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15969 (.I0(n1292), .I1(n1257), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15969.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15970 (.I0(n1290), .I1(n1255), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15970.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15971 (.I0(n1288), .I1(n1253), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15971.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15972 (.I0(n1286), .I1(n1251), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15972.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15973 (.I0(n1284), .I1(n1249), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15973.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15974 (.I0(n1282), .I1(n1247), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15974.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15975 (.I0(n1280), .I1(n1245), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15975.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15976 (.I0(n1278), .I1(n1243), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15976.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15977 (.I0(n1276), .I1(n1241), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15977.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15978 (.I0(n1274), .I1(n1239), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15978.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15979 (.I0(n1272), .I1(n1237), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15979.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15980 (.I0(n1266), .I1(n1235), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15980.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15981 (.I0(n1264), .I1(n1233), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15981.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15982 (.I0(n1263), .I1(n1232), .I2(n10511), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__15982.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__15983 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19] ), 
            .O(n10518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15983.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15984 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17] ), 
            .O(n10519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__15984.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__15985 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21] ), 
            .O(n10520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__15985.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__15986 (.I0(n10519), .I1(n10520), .I2(n10518), .I3(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11] ), 
            .O(n10521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__15986.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__15987 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12] ), 
            .I1(n10521), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__15987.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__15988 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9] ), 
            .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__15988.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__15989 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13] ), 
            .I1(n1922), .I2(n10521), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n343 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15989.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15990 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14] ), 
            .I1(n951), .I2(n10521), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15990.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15991 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15] ), 
            .I1(n948), .I2(n10521), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n341 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15991.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15992 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16] ), 
            .I1(n944), .I2(n10521), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15992.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15993 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17] ), 
            .I1(n942), .I2(n10521), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n339 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15993.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15994 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18] ), 
            .I1(n938), .I2(n10521), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15994.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15995 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19] ), 
            .I1(n936), .I2(n10521), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n337 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15995.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15996 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20] ), 
            .I1(n934), .I2(n10521), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15996.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__15997 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21] ), 
            .I1(n933), .I2(n10521), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__15997.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16001 (.I0(\u_axi4_ctrl/wframe_vsync_dly[3] ), .I1(\u_axi4_ctrl/wframe_vsync_dly[2] ), 
            .I2(\Axi0ResetReg[2] ), .O(\u_axi4_ctrl/n1469 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__16001.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__16002 (.I0(\u_axi4_ctrl/wframe_index[0] ), .I1(\u_axi4_ctrl/wframe_index[1] ), 
            .O(\u_axi4_ctrl/n317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16002.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16003 (.I0(\u_axi4_ctrl/wframe_vsync_dly[2] ), .I1(\u_axi4_ctrl/wframe_vsync_dly[3] ), 
            .O(\u_axi4_ctrl/equal_38/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__16003.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__16004 (.I0(\u_axi4_ctrl/wframe_index[0] ), .I1(\u_axi4_ctrl/wframe_index[1] ), 
            .O(\u_axi4_ctrl/n336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16004.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16005 (.I0(\u_axi4_ctrl/rframe_vsync_dly[2] ), .I1(\u_axi4_ctrl/rframe_vsync_dly[3] ), 
            .O(\u_axi4_ctrl/equal_47/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__16005.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__16006 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/rdata_cnt_dly[3] ), 
            .O(n10524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__16006.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__16007 (.I0(\u_axi4_ctrl/rdata_cnt_dly[4] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[5] ), 
            .I2(n10524), .O(n10525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__16007.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__16008 (.I0(DdrCtrl_RVALID_0), .I1(DdrCtrl_RREADY_0), .O(\u_axi4_ctrl/n379 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16008.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16009 (.I0(\u_axi4_ctrl/rdata_cnt_dly[6] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[7] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[8] ), .O(n10526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__16009.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__16010 (.I0(n10525), .I1(\u_axi4_ctrl/n379 ), .I2(n10526), 
            .O(\u_axi4_ctrl/n381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__16010.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__16011 (.I0(\u_axi4_ctrl/state[1] ), .I1(\u_axi4_ctrl/n381 ), 
            .I2(\u_axi4_ctrl/state[2] ), .O(n10527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__16011.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__16012 (.I0(DdrCtrl_BVALID_0), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(DdrCtrl_WREADY_0), .I3(DdrCtrl_WLAST_0), .O(n10528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__16012.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__16013 (.I0(n566), .I1(n567), .O(n10529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16013.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16014 (.I0(n431), .I1(n433), .I2(n435), .I3(n437), 
            .O(n10530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__16014.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__16015 (.I0(n439), .I1(n2526), .O(n10531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16015.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16016 (.I0(n10531), .I1(n10530), .I2(n429), .I3(n428), 
            .O(n10532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__16016.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__16017 (.I0(n10532), .I1(n10529), .I2(DdrCtrl_AREADY_0), 
            .I3(\u_axi4_ctrl/state[0] ), .O(n10533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__16017.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__16018 (.I0(n10533), .I1(n10528), .I2(\u_axi4_ctrl/state[2] ), 
            .I3(\u_axi4_ctrl/state[1] ), .O(n10534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__16018.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__16019 (.I0(\u_axi4_ctrl/state[0] ), .I1(DdrCtrl_AREADY_0), 
            .I2(n10527), .I3(n10534), .O(\u_axi4_ctrl/n389 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0 */ ;
    defparam LUT__16019.LUTMASK = 16'hffe0;
    EFX_LUT4 LUT__16020 (.I0(\u_axi4_ctrl/state[0] ), .I1(\u_axi4_ctrl/state[1] ), 
            .I2(\u_axi4_ctrl/state[2] ), .I3(n10529), .O(\u_axi4_ctrl/n405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__16020.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__16021 (.I0(\u_axi4_ctrl/state[0] ), .I1(\u_axi4_ctrl/state[1] ), 
            .I2(\u_axi4_ctrl/state[2] ), .I3(n10532), .O(n10535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__16021.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__16022 (.I0(n10535), .I1(\Axi0ResetReg[2] ), .O(\u_axi4_ctrl/n1476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__16022.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__16023 (.I0(DdrCtrl_WREADY_0), .I1(DdrCtrl_WVALID_0), .O(\u_axi4_ctrl/n363 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16023.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16024 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .O(\u_axi4_ctrl/n1544 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16024.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16029 (.I0(n662), .I1(n664), .I2(n666), .I3(n2355), 
            .O(n10536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__16029.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__16030 (.I0(n651), .I1(n652), .I2(n654), .I3(n656), 
            .O(n10537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__16030.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__16031 (.I0(n658), .I1(n660), .I2(n10536), .I3(n10537), 
            .O(n10538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__16031.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__16032 (.I0(\u_axi4_ctrl/n363 ), .I1(\u_axi4_ctrl/wfifo_empty ), 
            .I2(n10538), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__16032.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__16033 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
            .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .O(n10539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0990 */ ;
    defparam LUT__16033.LUTMASK = 16'h0990;
    EFX_LUT4 LUT__16034 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] ), 
            .I2(n10539), .O(n10540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__16034.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__16035 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .O(n10541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__16035.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__16036 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .O(n10542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__16036.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__16037 (.I0(n10541), .I1(n10542), .O(n10543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16037.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16038 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] ), .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), 
            .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .O(n10544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__16038.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__16039 (.I0(n10543), .I1(n10544), .I2(n10540), .I3(tvalid_o), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__16039.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__16040 (.I0(\u_axi4_ctrl/wframe_index[1] ), .I1(\u_axi4_ctrl/wframe_index[0] ), 
            .O(\u_axi4_ctrl/n316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16040.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16041 (.I0(\u_axi4_ctrl/n363 ), .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
            .O(ceg_net289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16041.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16042 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16042.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16043 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16043.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16044 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16044.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16045 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16045.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16046 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16046.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16047 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16047.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16048 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16048.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16049 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16049.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16050 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n7366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__16050.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__16051 (.I0(n5740), .I1(n7366), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16051.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16054 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] ), 
            .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .O(n10545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__16054.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__16055 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .O(n10546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__16055.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__16056 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .O(n10547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__16056.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__16057 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] ), 
            .O(n10548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__16057.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__16058 (.I0(n10546), .I1(n10547), .I2(n10548), .O(n10549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__16058.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__16059 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .I2(n10545), .I3(n10549), .O(n10550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__16059.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__16060 (.I0(lcd_de), .I1(\u_axi4_ctrl/rfifo_empty ), .I2(n10550), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__16060.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__16061 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12] ), 
            .O(n10551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0990 */ ;
    defparam LUT__16061.LUTMASK = 16'h0990;
    EFX_LUT4 LUT__16062 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .I2(n10551), .O(n10552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__16062.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__16063 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .O(n10553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__16063.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__16064 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] ), 
            .O(n10554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__16064.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__16065 (.I0(n10553), .I1(n10554), .O(n10555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16065.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16066 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] ), 
            .O(n10556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__16066.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__16067 (.I0(n10555), .I1(n10556), .I2(n10552), .I3(\u_axi4_ctrl/rfifo_wenb ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__16067.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__16068 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16068.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16069 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16069.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16070 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16070.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16071 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16071.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16072 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16072.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16073 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16073.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16074 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16074.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16075 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16075.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16076 (.I0(n5737), .I1(n5740), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16076.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16077 (.I0(n5734), .I1(n5737), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16077.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16078 (.I0(n5723), .I1(n5734), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16078.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16079 (.I0(n5660), .I1(n5723), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16079.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16080 (.I0(n5626), .I1(n5660), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16080.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16081 (.I0(n5623), .I1(n5626), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16081.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16082 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16082.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16083 (.I0(n5623), .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__16083.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__16084 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16084.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16085 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16085.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16086 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16086.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16087 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16087.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16088 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16088.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16089 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16089.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16090 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16090.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16091 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16091.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16092 (.I0(lcd_de), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
            .O(ceg_net296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16092.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16093 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16093.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16094 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF_frt_32_q ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16094.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16095 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16095.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16096 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16096.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16097 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16097.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16098 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16098.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16099 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16099.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16100 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16100.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16101 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16101.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16104 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16104.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16105 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[11] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16105.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16106 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16106.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16107 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16107.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16108 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16108.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16109 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16109.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16110 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16110.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16111 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16111.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16112 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .O(n10557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16112.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16113 (.I0(n10557), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__16113.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__16114 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .O(n10558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16114.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16115 (.I0(n10558), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__16115.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__16116 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .O(n10559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16116.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16117 (.I0(n10559), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__16117.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__16118 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .O(n10560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16118.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16119 (.I0(n10560), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__16119.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__16120 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .O(n10561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16120.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16121 (.I0(n10561), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__16121.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__16122 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] ), 
            .O(n10562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16122.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16123 (.I0(n10562), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__16123.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__16124 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] ), .I2(\u_axi4_ctrl/rfifo_empty ), 
            .O(n10563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16124.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16125 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] ), 
            .I2(\u_axi4_ctrl/rfifo_empty ), .I3(n10563), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h53ac */ ;
    defparam LUT__16125.LUTMASK = 16'h53ac;
    EFX_LUT4 LUT__16126 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] ), 
            .I2(\u_axi4_ctrl/rfifo_empty ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16126.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16127 (.I0(n10563), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16127.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16128 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16128.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16129 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16129.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16130 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16130.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16131 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16131.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16132 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16132.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16133 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16133.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16134 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16134.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16135 (.I0(\u_axi4_ctrl/wframe_index[0] ), .I1(\u_axi4_ctrl/wframe_index[1] ), 
            .O(\u_axi4_ctrl/n335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__16135.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__16136 (.I0(\u_axi4_ctrl/state[2] ), .I1(\u_axi4_ctrl/state[0] ), 
            .O(n10564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16136.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16137 (.I0(DdrCtrl_AREADY_0), .I1(DdrCtrl_BVALID_0), .I2(n10564), 
            .I3(\u_axi4_ctrl/state[1] ), .O(\u_axi4_ctrl/n1612 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3fa0 */ ;
    defparam LUT__16137.LUTMASK = 16'h3fa0;
    EFX_LUT4 LUT__16138 (.I0(\u_axi4_ctrl/state[2] ), .I1(\Axi0ResetReg[2] ), 
            .O(\u_axi4_ctrl/n1619 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__16138.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__16139 (.I0(n10527), .I1(n10535), .O(\u_axi4_ctrl/n387 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__16139.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__16140 (.I0(DdrCtrl_BVALID_0), .I1(DdrCtrl_BREADY_0), .O(\u_axi4_ctrl/n369 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16140.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16141 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .I1(n7838), .O(n7841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16141.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16142 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .I1(n7841), .O(n7844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16142.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16143 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .I1(n7850), .O(n7853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16143.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16144 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] ), 
            .I1(n7856), .O(n7859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16144.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16145 (.I0(\u_axi4_ctrl/rframe_vsync_dly[3] ), .I1(\u_axi4_ctrl/rframe_vsync_dly[2] ), 
            .I2(\Axi0ResetReg[2] ), .O(\u_axi4_ctrl/n1478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__16145.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__16146 (.I0(\u_axi4_ctrl/araddr[10] ), .I1(\u_axi4_ctrl/awaddr[10] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16146.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16147 (.I0(\u_axi4_ctrl/n405 ), .I1(\u_axi4_ctrl/n1476 ), 
            .O(ceg_net401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16147.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16148 (.I0(\u_axi4_ctrl/araddr[11] ), .I1(\u_axi4_ctrl/awaddr[11] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16148.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16149 (.I0(\u_axi4_ctrl/araddr[12] ), .I1(\u_axi4_ctrl/awaddr[12] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n695 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16149.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16150 (.I0(\u_axi4_ctrl/araddr[13] ), .I1(\u_axi4_ctrl/awaddr[13] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16150.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16151 (.I0(\u_axi4_ctrl/araddr[14] ), .I1(\u_axi4_ctrl/awaddr[14] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16151.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16152 (.I0(\u_axi4_ctrl/araddr[15] ), .I1(\u_axi4_ctrl/awaddr[15] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16152.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16153 (.I0(\u_axi4_ctrl/araddr[16] ), .I1(\u_axi4_ctrl/awaddr[16] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16153.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16154 (.I0(\u_axi4_ctrl/araddr[17] ), .I1(\u_axi4_ctrl/awaddr[17] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16154.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16155 (.I0(\u_axi4_ctrl/araddr[18] ), .I1(\u_axi4_ctrl/awaddr[18] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n689 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16155.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16156 (.I0(\u_axi4_ctrl/araddr[19] ), .I1(\u_axi4_ctrl/awaddr[19] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n688 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16156.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16157 (.I0(\u_axi4_ctrl/araddr[20] ), .I1(\u_axi4_ctrl/awaddr[20] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n687 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16157.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16158 (.I0(\u_axi4_ctrl/araddr[21] ), .I1(\u_axi4_ctrl/awaddr[21] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n686 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16158.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16159 (.I0(\u_axi4_ctrl/araddr[22] ), .I1(\u_axi4_ctrl/awaddr[22] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n685 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16159.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16160 (.I0(\u_axi4_ctrl/araddr[23] ), .I1(\u_axi4_ctrl/awaddr[23] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16160.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16161 (.I0(\u_axi4_ctrl/rframe_index[0] ), .I1(\u_axi4_ctrl/wframe_index[0] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n683 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16161.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16162 (.I0(\u_axi4_ctrl/rframe_index[1] ), .I1(\u_axi4_ctrl/wframe_index[1] ), 
            .I2(n10535), .O(\u_axi4_ctrl/n682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__16162.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__16163 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .O(\u_axi4_ctrl/n1499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16163.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16164 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .O(\u_axi4_ctrl/n1504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__16164.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__16165 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/wdata_cnt_dly[3] ), 
            .O(\u_axi4_ctrl/n1509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__16165.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__16166 (.I0(\u_axi4_ctrl/wdata_cnt_dly[4] ), .I1(n10069), 
            .O(\u_axi4_ctrl/n1514 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16166.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16167 (.I0(\u_axi4_ctrl/wdata_cnt_dly[4] ), .I1(n10069), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[5] ), .O(\u_axi4_ctrl/n1519 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__16167.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__16168 (.I0(\u_axi4_ctrl/wdata_cnt_dly[6] ), .I1(n10070), 
            .O(\u_axi4_ctrl/n1524 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16168.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16169 (.I0(\u_axi4_ctrl/wdata_cnt_dly[6] ), .I1(n10070), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[7] ), .O(\u_axi4_ctrl/n1529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__16169.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__16170 (.I0(\u_axi4_ctrl/wdata_cnt_dly[6] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[7] ), 
            .I2(n10070), .I3(\u_axi4_ctrl/wdata_cnt_dly[8] ), .O(\u_axi4_ctrl/n1534 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__16170.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__16171 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[2] ), .O(\u_axi4_ctrl/n1549 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__16171.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__16172 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/rdata_cnt_dly[3] ), 
            .O(\u_axi4_ctrl/n1554 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__16172.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__16173 (.I0(\u_axi4_ctrl/rdata_cnt_dly[4] ), .I1(n10524), 
            .O(\u_axi4_ctrl/n1559 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16173.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16174 (.I0(\u_axi4_ctrl/rdata_cnt_dly[4] ), .I1(n10524), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[5] ), .O(\u_axi4_ctrl/n1564 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__16174.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__16175 (.I0(\u_axi4_ctrl/rdata_cnt_dly[6] ), .I1(n10525), 
            .O(\u_axi4_ctrl/n1569 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16175.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16176 (.I0(\u_axi4_ctrl/rdata_cnt_dly[6] ), .I1(n10525), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[7] ), .O(\u_axi4_ctrl/n1574 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__16176.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__16177 (.I0(\u_axi4_ctrl/rdata_cnt_dly[6] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[7] ), 
            .I2(n10525), .I3(\u_axi4_ctrl/rdata_cnt_dly[8] ), .O(\u_axi4_ctrl/n1579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__16177.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__16178 (.I0(\u_lcd_driver/vcnt[3] ), .I1(\u_lcd_driver/vcnt[4] ), 
            .I2(\u_lcd_driver/vcnt[5] ), .I3(\u_lcd_driver/vcnt[6] ), .O(n10565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__16178.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__16179 (.I0(\u_lcd_driver/n76 ), .I1(\u_lcd_driver/n75 ), 
            .O(n10566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16179.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16180 (.I0(\u_lcd_driver/vcnt[2] ), .I1(\u_lcd_driver/vcnt[1] ), 
            .I2(n10565), .I3(\u_lcd_driver/vcnt[7]~FF_frt_39_q ), .O(n10567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__16180.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__16181 (.I0(n10567), .I1(\u_lcd_driver/vcnt[9] ), .I2(\u_lcd_driver/vcnt[11] ), 
            .I3(\u_lcd_driver/vcnt[10] ), .O(n10568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__16181.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__16182 (.I0(\u_lcd_driver/vcnt[0] ), .I1(n10568), .O(\u_lcd_driver/n83 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16182.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16183 (.I0(\u_lcd_driver/hcnt[0] ), .I1(\u_lcd_driver/hcnt[1] ), 
            .I2(\u_lcd_driver/hcnt[2] ), .I3(\u_lcd_driver/hcnt[3] ), .O(n10569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__16183.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__16184 (.I0(\u_lcd_driver/hcnt[4] ), .I1(\u_lcd_driver/hcnt[5] ), 
            .I2(n10569), .O(n10570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__16184.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__16185 (.I0(\u_lcd_driver/hcnt[6] ), .I1(\u_lcd_driver/hcnt[7] ), 
            .I2(\u_lcd_driver/hcnt[9] ), .I3(\u_lcd_driver/hcnt[11] ), .O(n10571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__16185.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__16186 (.I0(\u_lcd_driver/hcnt[8] ), .I1(\u_lcd_driver/hcnt[10] ), 
            .I2(n10570), .I3(n10571), .O(\u_lcd_driver/equal_17/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__16186.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__16187 (.I0(\u_lcd_driver/hcnt[4] ), .I1(\u_lcd_driver/hcnt[3] ), 
            .I2(\u_lcd_driver/hcnt[5] ), .O(n10572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__16187.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__16188 (.I0(\u_lcd_driver/hcnt[8] ), .I1(\u_lcd_driver/hcnt[10] ), 
            .I2(n10572), .I3(n10571), .O(\u_lcd_driver/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__16188.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__16189 (.I0(\u_lcd_driver/n82 ), .I1(\u_lcd_driver/n83 ), 
            .I2(\u_lcd_driver/n79 ), .I3(\u_lcd_driver/n78 ), .O(n10573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__16189.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__16190 (.I0(\u_lcd_driver/n81 ), .I1(\u_lcd_driver/n80 ), 
            .I2(n10573), .O(n10574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__16190.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__16191 (.I0(\u_lcd_driver/vcnt[6] ), .I1(\u_lcd_driver/vcnt[9] ), 
            .I2(\u_lcd_driver/vcnt[7]~FF_frt_39_q ), .O(n10575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__16191.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__16192 (.I0(\u_lcd_driver/vcnt[10] ), .I1(\u_lcd_driver/vcnt[11] ), 
            .I2(\u_lcd_driver/vcnt[2]~FF_frt_40_q ), .I3(n10575), .O(\u_lcd_driver/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__16192.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__16193 (.I0(\u_lcd_driver/vcnt[0] ), .I1(\u_lcd_driver/vcnt[1] ), 
            .I2(\u_lcd_driver/vcnt[2] ), .O(n10576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__16193.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__16194 (.I0(\u_lcd_driver/vcnt[3] ), .I1(n10576), .I2(\u_lcd_driver/vcnt[4] ), 
            .I3(\u_lcd_driver/vcnt[5] ), .O(n10577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h07e0 */ ;
    defparam LUT__16194.LUTMASK = 16'h07e0;
    EFX_LUT4 LUT__16195 (.I0(n10575), .I1(\u_lcd_driver/vcnt[6] ), .I2(n10577), 
            .I3(\u_lcd_driver/vcnt[5] ), .O(n10578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__16195.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__16196 (.I0(\u_lcd_driver/vcnt[7]~FF_frt_39_q ), .I1(\u_lcd_driver/vcnt[5] ), 
            .I2(n10578), .I3(\u_lcd_driver/vcnt[9] ), .O(n10579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf530 */ ;
    defparam LUT__16196.LUTMASK = 16'hf530;
    EFX_LUT4 LUT__16197 (.I0(\u_lcd_driver/n28 ), .I1(\u_lcd_driver/n29 ), 
            .I2(\u_lcd_driver/n27 ), .O(n10580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__16197.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__16198 (.I0(\u_lcd_driver/n26 ), .I1(\u_lcd_driver/n25 ), 
            .I2(n10580), .I3(\u_lcd_driver/n24 ), .O(n10581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h01fe */ ;
    defparam LUT__16198.LUTMASK = 16'h01fe;
    EFX_LUT4 LUT__16199 (.I0(\u_lcd_driver/vcnt[10] ), .I1(\u_lcd_driver/vcnt[11] ), 
            .I2(\u_lcd_driver/hcnt[11] ), .I3(\u_lcd_driver/hcnt[8]~FF_frt_41_q ), 
            .O(n10582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__16199.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__16200 (.I0(n10579), .I1(n10582), .O(\u_lcd_driver/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16200.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16201 (.I0(\u_lcd_driver/vcnt[2]~FF_frt_40_q ), .I1(\u_lcd_driver/vcnt[6] ), 
            .I2(\u_lcd_driver/vcnt[7]~FF_frt_39_q ), .O(n10583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__16201.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__16202 (.I0(\u_lcd_driver/vcnt[9] ), .I1(n10583), .I2(n10582), 
            .O(\u_lcd_driver/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__16202.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__16203 (.I0(\u_lcd_driver/hcnt[9] ), .I1(\u_lcd_driver/hcnt[8] ), 
            .I2(\u_lcd_driver/hcnt[10] ), .I3(\u_lcd_driver/hcnt[11] ), 
            .O(n10584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__16203.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__16204 (.I0(n10571), .I1(n10570), .I2(n10584), .O(n10585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__16204.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__16205 (.I0(\u_lcd_driver/hcnt[0] ), .I1(n10585), .O(\u_lcd_driver/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__16205.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__16206 (.I0(n3039), .I1(n10568), .O(\u_lcd_driver/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16206.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16207 (.I0(n407), .I1(n10568), .O(\u_lcd_driver/n81 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16207.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16208 (.I0(n405), .I1(n10568), .O(\u_lcd_driver/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16208.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16209 (.I0(n403), .I1(n10568), .O(\u_lcd_driver/n79 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16209.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16210 (.I0(n401), .I1(n10568), .O(\u_lcd_driver/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16210.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16211 (.I0(n399), .I1(n10568), .O(\u_lcd_driver/n77 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16211.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16212 (.I0(n397), .I1(n10568), .O(\u_lcd_driver/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16212.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16213 (.I0(n395), .I1(n10568), .O(\u_lcd_driver/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16213.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16214 (.I0(n393), .I1(n10568), .O(\u_lcd_driver/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16214.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16215 (.I0(n391), .I1(n10568), .O(\u_lcd_driver/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16215.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16216 (.I0(n390), .I1(n10568), .O(\u_lcd_driver/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__16216.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__16217 (.I0(n10585), .I1(n2543), .O(\u_lcd_driver/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16217.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16218 (.I0(n10585), .I1(n426), .O(\u_lcd_driver/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16218.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16219 (.I0(n10585), .I1(n424), .O(\u_lcd_driver/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16219.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16220 (.I0(n10585), .I1(n422), .O(\u_lcd_driver/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16220.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16221 (.I0(n10585), .I1(n420), .O(\u_lcd_driver/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16221.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16222 (.I0(n10585), .I1(n418), .O(\u_lcd_driver/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16222.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16223 (.I0(n10585), .I1(n416), .O(\u_lcd_driver/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16223.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16224 (.I0(n10585), .I1(n414), .O(\u_lcd_driver/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16224.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16225 (.I0(n10585), .I1(n412), .O(\u_lcd_driver/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16225.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16226 (.I0(n10585), .I1(n410), .O(\u_lcd_driver/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16226.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16227 (.I0(n10585), .I1(n409), .O(\u_lcd_driver/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__16227.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__16228 (.I0(n10322), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .I2(n10297), .I3(\u_rgb2dvi/enc_0/acc[4] ), .O(n10586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3c27 */ ;
    defparam LUT__16228.LUTMASK = 16'h3c27;
    EFX_LUT4 LUT__16229 (.I0(\u_rgb2dvi/enc_0/acc[4] ), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .I2(n10323), .I3(n10586), .O(n10587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88c7 */ ;
    defparam LUT__16229.LUTMASK = 16'h88c7;
    EFX_LUT4 LUT__16230 (.I0(lcd_hs), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q ), 
            .I2(n10587), .I3(lcd_de), .O(\u_rgb2dvi/enc_0/n866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3aa */ ;
    defparam LUT__16230.LUTMASK = 16'hc3aa;
    EFX_LUT4 LUT__16231 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_24_q ), .O(n10588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__16231.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__16232 (.I0(lcd_hs), .I1(n10587), .I2(n10588), .I3(lcd_de), 
            .O(\u_rgb2dvi/enc_0/n768 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3aa */ ;
    defparam LUT__16232.LUTMASK = 16'hc3aa;
    EFX_LUT4 LUT__16233 (.I0(lcd_hs), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_q ), 
            .I2(n10587), .I3(lcd_de), .O(\u_rgb2dvi/enc_0/n774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__16233.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__16234 (.I0(\u_lcd_driver/r_lcd_dv ), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_11_q ), 
            .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), .O(n10589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7c7c */ ;
    defparam LUT__16234.LUTMASK = 16'h7c7c;
    EFX_LUT4 LUT__16235 (.I0(lcd_hs), .I1(n10587), .I2(n10589), .I3(lcd_de), 
            .O(\u_rgb2dvi/enc_0/n780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__16235.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__16236 (.I0(lcd_hs), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_q ), 
            .I2(n10587), .I3(lcd_de), .O(\u_rgb2dvi/enc_0/n786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__16236.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__16237 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26_q ), .O(n10590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16237.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16238 (.I0(lcd_hs), .I1(n10587), .I2(n10590), .I3(lcd_de), 
            .O(\u_rgb2dvi/enc_0/n792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3aa */ ;
    defparam LUT__16238.LUTMASK = 16'hc3aa;
    EFX_LUT4 LUT__16239 (.I0(lcd_hs), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27_q ), 
            .I2(n10587), .I3(lcd_de), .O(\u_rgb2dvi/enc_0/n798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__16239.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__16240 (.I0(lcd_hs), .I1(n10319), .I2(n10587), .I3(lcd_de), 
            .O(\u_rgb2dvi/enc_0/n804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3aa */ ;
    defparam LUT__16240.LUTMASK = 16'hc3aa;
    EFX_LUT4 LUT__16241 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .I1(lcd_hs), .I2(lcd_de), .O(\u_rgb2dvi/enc_0/n810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__16241.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__16242 (.I0(n10587), .I1(lcd_vs), .I2(lcd_hs), .I3(lcd_de), 
            .O(\u_rgb2dvi/enc_0/n816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h55c3 */ ;
    defparam LUT__16242.LUTMASK = 16'h55c3;
    EFX_LUT4 LUT__16243 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .I1(n10312), .I2(n10315), .I3(n10297), .O(\u_rgb2dvi/enc_1/q_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h35cd */ ;
    defparam LUT__16243.LUTMASK = 16'h35cd;
    EFX_LUT4 LUT__16244 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q ), .I1(\u_rgb2dvi/enc_1/q_out[9] ), 
            .O(\u_rgb2dvi/enc_1/q_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16244.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16245 (.I0(n10588), .I1(\u_rgb2dvi/enc_1/q_out[9] ), .O(\u_rgb2dvi/enc_1/q_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16245.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16246 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_q ), .I1(\u_rgb2dvi/enc_1/q_out[9] ), 
            .O(\u_rgb2dvi/enc_1/q_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16246.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16247 (.I0(n10589), .I1(\u_rgb2dvi/enc_1/q_out[9] ), .O(\u_rgb2dvi/enc_1/q_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__16247.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__16248 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_q ), 
            .I1(\u_rgb2dvi/enc_1/q_out[9] ), .O(\u_rgb2dvi/enc_1/q_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16248.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16249 (.I0(n10590), .I1(\u_rgb2dvi/enc_1/q_out[9] ), .O(\u_rgb2dvi/enc_1/q_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16249.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16250 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27_q ), 
            .I1(\u_rgb2dvi/enc_1/q_out[9] ), .O(\u_rgb2dvi/enc_1/q_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16250.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16251 (.I0(n10319), .I1(\u_rgb2dvi/enc_1/q_out[9] ), .O(\u_rgb2dvi/enc_1/q_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16251.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16252 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q ), 
            .I1(n10299), .I2(n10304), .I3(n10297), .O(\u_rgb2dvi/enc_2/q_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h35cd */ ;
    defparam LUT__16252.LUTMASK = 16'h35cd;
    EFX_LUT4 LUT__16253 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q ), .I1(\u_rgb2dvi/enc_2/q_out[9] ), 
            .O(\u_rgb2dvi/enc_2/q_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16253.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16254 (.I0(n10588), .I1(\u_rgb2dvi/enc_2/q_out[9] ), .O(\u_rgb2dvi/enc_2/q_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16254.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16255 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_q ), .I1(\u_rgb2dvi/enc_2/q_out[9] ), 
            .O(\u_rgb2dvi/enc_2/q_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16255.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16256 (.I0(n10589), .I1(\u_rgb2dvi/enc_2/q_out[9] ), .O(\u_rgb2dvi/enc_2/q_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__16256.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__16257 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_q ), 
            .I1(\u_rgb2dvi/enc_2/q_out[9] ), .O(\u_rgb2dvi/enc_2/q_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16257.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16258 (.I0(n10590), .I1(\u_rgb2dvi/enc_2/q_out[9] ), .O(\u_rgb2dvi/enc_2/q_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16258.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16259 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27_q ), 
            .I1(\u_rgb2dvi/enc_2/q_out[9] ), .O(\u_rgb2dvi/enc_2/q_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16259.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16260 (.I0(n10319), .I1(\u_rgb2dvi/enc_2/q_out[9] ), .O(\u_rgb2dvi/enc_2/q_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__16260.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__16261 (.I0(\r_hdmi_tx0_o[6] ), .I1(\w_hdmi_txd0[1] ), 
            .I2(rc_hdmi_tx), .O(n591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16261.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16262 (.I0(\r_hdmi_tx0_o[7] ), .I1(\w_hdmi_txd0[2] ), 
            .I2(rc_hdmi_tx), .O(n590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__16262.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__16263 (.I0(\r_hdmi_tx0_o[8] ), .I1(\w_hdmi_txd0[3] ), 
            .I2(rc_hdmi_tx), .O(n589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16263.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16264 (.I0(\r_hdmi_tx0_o[9] ), .I1(\w_hdmi_txd0[4] ), 
            .I2(rc_hdmi_tx), .O(n588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__16264.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__16265 (.I0(\r_hdmi_tx1_o[6] ), .I1(\w_hdmi_txd1[1] ), 
            .I2(rc_hdmi_tx), .O(n602_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16265.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16266 (.I0(\r_hdmi_tx1_o[7] ), .I1(\w_hdmi_txd1[2] ), 
            .I2(rc_hdmi_tx), .O(n601_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__16266.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__16267 (.I0(\r_hdmi_tx1_o[8] ), .I1(\w_hdmi_txd1[3] ), 
            .I2(rc_hdmi_tx), .O(n600_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16267.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16268 (.I0(\r_hdmi_tx1_o[9] ), .I1(\w_hdmi_txd1[4] ), 
            .I2(rc_hdmi_tx), .O(n599_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__16268.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__16269 (.I0(\r_hdmi_tx2_o[6] ), .I1(\w_hdmi_txd2[1] ), 
            .I2(rc_hdmi_tx), .O(n613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16269.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16270 (.I0(\r_hdmi_tx2_o[7] ), .I1(\w_hdmi_txd2[2] ), 
            .I2(rc_hdmi_tx), .O(n612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__16270.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__16271 (.I0(\r_hdmi_tx1_o[8] ), .I1(\w_hdmi_txd2[3] ), 
            .I2(rc_hdmi_tx), .O(n611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__16271.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__16272 (.I0(\r_hdmi_tx2_o[9] ), .I1(\w_hdmi_txd2[4] ), 
            .I2(rc_hdmi_tx), .O(n610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__16272.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__16357 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
            .O(DdrCtrl_CFG_SEQ_RST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16357.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16381 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[0] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16381.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16382 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[1] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16382.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16383 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[2] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16383.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16384 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[3] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16384.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16385 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[4] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16385.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16386 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[5] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16386.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16387 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[6] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16387.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16388 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[7] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16388.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16389 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[8] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16389.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16390 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[9] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16390.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16391 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16391.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16392 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16392.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16394 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[0] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16394.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16395 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[1] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16395.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16396 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[2] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16396.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16397 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[3] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16397.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16398 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[4] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16398.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16399 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[5] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16399.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16400 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[6] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16400.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16401 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[7] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16401.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16402 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[8] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16402.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16403 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[9] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16403.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16404 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16404.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16405 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16405.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16406 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[8] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16406.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16407 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[9] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16407.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16408 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16408.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16409 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16409.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16410 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[8] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16410.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16411 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[9] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16411.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16412 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16412.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__16413 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__16413.LUTMASK = 16'h5555;
    EFX_LUT4 \u_lcd_driver/vcnt[2]~FF_frt_40_rtinv  (.I0(\u_lcd_driver/vcnt[2]~FF_frt_40_q_pinv ), 
            .O(\u_lcd_driver/vcnt[2]~FF_frt_40_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \u_lcd_driver/vcnt[2]~FF_frt_40_rtinv .LUTMASK = 16'h5555;
    EFX_LUT4 \u_lcd_driver/vcnt[7]~FF_frt_39_rtinv  (.I0(\u_lcd_driver/vcnt[7]~FF_frt_39_q_pinv ), 
            .O(\u_lcd_driver/vcnt[7]~FF_frt_39_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \u_lcd_driver/vcnt[7]~FF_frt_39_rtinv .LUTMASK = 16'h5555;
    EFX_FF \u_lcd_driver/hcnt[8]~FF_frt_41  (.D(n10581), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[8]~FF_frt_41_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[8]~FF_frt_41 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF_frt_41 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF_frt_41 .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF_frt_41 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF_frt_41 .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF_frt_41 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF_frt_41 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[2]~FF_frt_40  (.D(n10574), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[2]~FF_frt_40_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[2]~FF_frt_40 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[2]~FF_frt_40 .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF_frt_40 .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF_frt_40 .D_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF_frt_40 .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF_frt_40 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF_frt_40 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38  (.D(n10302), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_frt_38 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_rtinv  (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q_pinv ), 
            .O(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q )) /* verific LUTMASK=16'h5555, EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_rtinv .LUTMASK = 16'h5555;
    EFX_FF \u_lcd_driver/vcnt[7]~FF_frt_39  (.D(n10566), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[7]~FF_frt_39_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[7]~FF_frt_39 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[7]~FF_frt_39 .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF_frt_39 .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF_frt_39 .D_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF_frt_39 .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF_frt_39 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF_frt_39 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28  (.D(n8411), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_28_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_28 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26  (.D(n10291), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_20_frt_26 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27  (.D(n10295), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_frt_27 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25  (.D(n8110), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25_q_pinv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25 .D_POLARITY = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_16_frt_21_frt_25 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_11  (.D(n10266), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_11_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_11 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_11 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_11 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_11 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_11 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_11 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_11 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10  (.D(n10272), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_24  (.D(n10293), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_24_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_24 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_24 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_24 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_24 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_24 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_24 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_24 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_dv~FF_frt_7  (.D(n10269), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\u_lcd_driver/r_lcd_dv~FF_frt_7_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22  (.D(n10284), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_10_frt_22 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0  (.D(n7826), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true", INIT_VALUE=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .SR_SYNC_PRIORITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_8d8d6396_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_8d8d6396_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_8d8d6396_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_8d8d6396_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_8d8d6396_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_8d8d6396_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_16_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_16_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_16_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_16_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_16_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_16_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_16_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_16_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__16_1_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__16_1_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__16_1_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__16_1_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__16_1_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__16_1_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__16_1_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__16_1_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_8d8d6396__1_1_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_MULT_8d8d6396_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_MULT_8d8d6396_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_MULT_8d8d6396_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_MULT_8d8d6396_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_214
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_215
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_216
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_217
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_218
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_219
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_220
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_221
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_222
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_223
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_224
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_225
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_226
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_227
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_228
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_229
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_230
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_231
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_232
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_233
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_234
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_235
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_236
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_237
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_238
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_239
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_240
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_241
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_242
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_243
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_244
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_245
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_246
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_247
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_248
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_249
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_250
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_251
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_252
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_253
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_254
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_255
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_256
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_257
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_258
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_259
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_260
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_261
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_262
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_263
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_264
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_265
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_266
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_267
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_268
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_269
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_270
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_271
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_272
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_273
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_274
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_275
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_276
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_277
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_278
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_279
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_280
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_281
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_282
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_283
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_284
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_285
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_286
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_287
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_288
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_289
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_290
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_291
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_292
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_293
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_294
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_295
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_296
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_8d8d6396_297
// module not written out since it is a black box. 
//



//
// Verific Verilog Description of module T35_Sensor_DDR3_LCD_Test
//

module T35_Sensor_DDR3_LCD_Test (Axi_Clk, tx_slowclk, tx_fastclk, pll_clk_200m, 
            hdmi_clk1x_i, hdmi_clk2x_i, hdmi_clk5x_i, PllLocked, DdrCtrl_CFG_RST_N, 
            DdrCtrl_CFG_SEQ_RST, DdrCtrl_CFG_SEQ_START, DdrCtrl_AID_0, 
            DdrCtrl_AADDR_0, DdrCtrl_ALEN_0, DdrCtrl_ASIZE_0, DdrCtrl_ABURST_0, 
            DdrCtrl_ALOCK_0, DdrCtrl_AVALID_0, DdrCtrl_AREADY_0, DdrCtrl_ATYPE_0, 
            DdrCtrl_WID_0, DdrCtrl_WDATA_0, DdrCtrl_WSTRB_0, DdrCtrl_WLAST_0, 
            DdrCtrl_WVALID_0, DdrCtrl_WREADY_0, DdrCtrl_RID_0, DdrCtrl_RDATA_0, 
            DdrCtrl_RLAST_0, DdrCtrl_RVALID_0, DdrCtrl_RREADY_0, DdrCtrl_RRESP_0, 
            DdrCtrl_BID_0, DdrCtrl_BVALID_0, DdrCtrl_BREADY_0, LED, 
            cmos_sclk, cmos_sdat_IN, cmos_sdat_OUT, cmos_sdat_OE, cmos_pclk, 
            cmos_vsync, cmos_href, cmos_data, cmos_ctl0, cmos_ctl1, 
            cmos_ctl2, cmos_ctl3, hdmi_tx0_o, hdmi_tx1_o, hdmi_tx2_o, 
            hdmi_txc_o, lcd_pwm, lvds_tx_clk_DATA, lvds_tx0_DATA, lvds_tx1_DATA, 
            lvds_tx2_DATA, lvds_tx3_DATA);
    input Axi_Clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input tx_slowclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input tx_fastclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input pll_clk_200m /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input hdmi_clk1x_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input hdmi_clk2x_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input hdmi_clk5x_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [1:0]PllLocked /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_CFG_RST_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_CFG_SEQ_RST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_CFG_SEQ_START /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_AID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [31:0]DdrCtrl_AADDR_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_ALEN_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [2:0]DdrCtrl_ASIZE_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]DdrCtrl_ABURST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]DdrCtrl_ALOCK_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_AVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input DdrCtrl_AREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_ATYPE_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_WID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [127:0]DdrCtrl_WDATA_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [15:0]DdrCtrl_WSTRB_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_WLAST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_WVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input DdrCtrl_WREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]DdrCtrl_RID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [127:0]DdrCtrl_RDATA_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_RLAST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_RVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_RREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [1:0]DdrCtrl_RRESP_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]DdrCtrl_BID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_BVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_BREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]LED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output cmos_sclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input cmos_sdat_IN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output cmos_sdat_OUT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output cmos_sdat_OE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input cmos_pclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input cmos_vsync /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input cmos_href /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]cmos_data /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output cmos_ctl0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input cmos_ctl1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output cmos_ctl2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output cmos_ctl3 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_tx0_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_tx1_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_tx2_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [4:0]hdmi_txc_o /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output lcd_pwm /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx_clk_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx0_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx1_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx2_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx3_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    wire \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire n2105_2;
    wire n592_2;
    wire n603_2;
    wire n614_2;
    wire n9_2;
    wire n2091_2;
    wire \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]  /* verific async_reg="true" */ ;
    wire \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]  /* verific async_reg="true" */ ;
    wire n197_2;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire n602_2;
    wire n601_2;
    
    wire n176, n177, \ResetShiftReg[0] , \Axi0ResetReg[0] , r_hdmi_rst_n, 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n98 , rc_hdmi_tx, \PowerOnResetCnt[0] , 
        \ResetShiftReg[1] , \Axi0ResetReg[1] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] , n197, n198, \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] , n219, n220, \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] , 
        n222, n223, \u_i2c_timing_ctrl_16reg_16bit/current_state[1] , 
        \u_i2c_timing_ctrl_16reg_16bit/current_state[0] , \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en , \i2c_config_index[0] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3] , \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2] , 
        \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1] , \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0] , \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5 , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4 , \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3 , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2 , \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1 , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_ack , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0] , \u_i2c_timing_ctrl_16reg_16bit/current_state[2] , 
        \u_i2c_timing_ctrl_16reg_16bit/current_state[3] , \u_i2c_timing_ctrl_16reg_16bit/current_state[4] , 
        \i2c_config_index[1] , \i2c_config_index[2] , \i2c_config_index[3] , 
        \i2c_config_index[4] , \i2c_config_index[5] , \i2c_config_index[6] , 
        \i2c_config_index[7] , \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] , \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] , \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3] , \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5] , \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17] , \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18] , 
        \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19] , n336, n337, n338, 
        n339, n340, n341, n342, n343, n344, n345, n346, n347, 
        n348, n349, n350, n351, n352, n353, n354, n355, n356, 
        n357, n358, n359, n360, n361, n362, n363, n364, n365, 
        n366, n367, n368, n369, n370, n371, n372, n373, n374, 
        n375, n376, n377, n378, n379, n380, n381, n382, n383, 
        n384, n385, n386, n387, n388, n389, n390, n391, n392, 
        n393, n394, n395, n396, n397, n398, n399, n400, n401, 
        n402, n403, n404, n405, n406, n407, n408, n409, n410, 
        n411, n412, n413, n414, n415, n416, n417, n418, n419, 
        n420, n421, n422, n423, n424, n425, n426, n427, n428, 
        n429, n430, n431, \u_CMOS_Capture_RAW_Gray/cmos_href_r[0] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0] , \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5] , n443, n444, \u_CMOS_Capture_RAW_Gray/line_cnt[0] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4] , \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7] , \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3] , n457, \u_CMOS_Capture_RAW_Gray/frame_sync_flag , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5] , \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2] , \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3] , 
        n464, n465, n466, n467, \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2] , 
        \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1] , \u_CMOS_Capture_RAW_Gray/cmos_href_r[1] , 
        n479, n480, \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] , \u_CMOS_Capture_RAW_Gray/line_cnt[1] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[2] , \u_CMOS_Capture_RAW_Gray/line_cnt[3] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[4] , \u_CMOS_Capture_RAW_Gray/line_cnt[5] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[6] , \u_CMOS_Capture_RAW_Gray/line_cnt[7] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[8] , \u_CMOS_Capture_RAW_Gray/line_cnt[9] , 
        \u_CMOS_Capture_RAW_Gray/line_cnt[10] , \u_CMOS_Capture_RAW_Gray/line_cnt[11] , 
        \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] , n524, n525, n534, 
        n535, n536, n537, n538, n539, n540, n541, n542, n543, 
        n544, n545, n546, n547, n548, n549, n550, n551, n552, 
        n553, n554, n555, n556, n557, n558, n559, n561, \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1] , 
        n575, n576, \u_sensor_frame_count/delay_cnt[9] , \u_sensor_frame_count/delay_cnt[8] , 
        \u_sensor_frame_count/delay_cnt[7] , \u_sensor_frame_count/delay_cnt[6] , 
        n597, \u_sensor_frame_count/delay_cnt[5] , \u_sensor_frame_count/delay_cnt[4] , 
        \u_sensor_frame_count/delay_cnt[1] , n601, n602, \u_sensor_frame_count/cmos_fps_cnt[0] , 
        \u_sensor_frame_count/delay_cnt[3] , \u_sensor_frame_count/delay_cnt[2] , 
        \u_sensor_frame_count/delay_cnt[0] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n105 , 
        \u_sensor_frame_count/cmos_vsync_r[0] , \u_sensor_frame_count/delay_cnt[10] , 
        \u_sensor_frame_count/delay_cnt[11] , \u_sensor_frame_count/delay_cnt[12] , 
        \u_sensor_frame_count/delay_cnt[13] , \u_sensor_frame_count/delay_cnt[14] , 
        \u_sensor_frame_count/delay_cnt[15] , \u_sensor_frame_count/delay_cnt[16] , 
        \u_sensor_frame_count/delay_cnt[17] , \u_sensor_frame_count/delay_cnt[18] , 
        \u_sensor_frame_count/delay_cnt[19] , \u_sensor_frame_count/delay_cnt[20] , 
        \u_sensor_frame_count/delay_cnt[21] , \u_sensor_frame_count/delay_cnt[22] , 
        \u_sensor_frame_count/delay_cnt[23] , \u_sensor_frame_count/delay_cnt[24] , 
        \u_sensor_frame_count/delay_cnt[25] , \u_sensor_frame_count/delay_cnt[26] , 
        \u_sensor_frame_count/delay_cnt[27] , n629, \u_sensor_frame_count/cmos_fps_cnt[2] , 
        \u_sensor_frame_count/cmos_fps_cnt[3] , \u_sensor_frame_count/cmos_fps_cnt[4] , 
        \u_sensor_frame_count/cmos_fps_cnt[5] , \u_sensor_frame_count/cmos_fps_cnt[6] , 
        \u_sensor_frame_count/cmos_fps_cnt[7] , \u_sensor_frame_count/cmos_fps_cnt[8] , 
        n639, n641, n642, n643, n644, n645, n646, n647, n648, 
        n649, n650, n651, n652, n653, n654, n655, n656, n657, 
        n658, n659, n660, n661, n662, n663, n664, n665, n666, 
        n667, n668, n669, n670, n671, n672, \u_sensor_frame_count/cmos_vsync_r[1] , 
        n681, n682, n683, n684, \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n99 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n102 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n104 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n96 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n93 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n90 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n87 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n84 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n101 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n95 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n92 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n89 , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n86 , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n83 , 
        n703, n704, \u_afifo_buf/u_efx_fifo_top/waddr[9] , \u_afifo_buf/u_efx_fifo_top/waddr[8] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[0] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[1] , empty, \u_afifo_buf/u_efx_fifo_top/waddr[6] , 
        n712, n713, \u_afifo_buf/u_efx_fifo_top/waddr[5] , n715, n716, 
        \u_afifo_buf/u_efx_fifo_top/raddr[0] , n718, n719, \u_afifo_buf/u_efx_fifo_top/waddr[4] , 
        n721, n722, n723, n724, \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[3] , \u_afifo_buf/u_efx_fifo_top/waddr[2] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[11] , 
        \u_afifo_buf/u_efx_fifo_top/waddr[12] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] , 
        n735, n736, n737, n738, n739, n740, n741, n742, n743, 
        n744, n745, n746, n747, n748, n749, n750, n751, n752, 
        n753, n754, n755, \u_afifo_buf/u_efx_fifo_top/raddr[1] , \u_afifo_buf/u_efx_fifo_top/raddr[2] , 
        \u_afifo_buf/u_efx_fifo_top/raddr[3] , \u_afifo_buf/u_efx_fifo_top/raddr[4] , 
        \u_afifo_buf/u_efx_fifo_top/raddr[5] , \u_afifo_buf/u_efx_fifo_top/raddr[6] , 
        \u_afifo_buf/u_efx_fifo_top/raddr[7] , \u_afifo_buf/u_efx_fifo_top/raddr[8] , 
        \u_afifo_buf/u_efx_fifo_top/raddr[9] , \u_afifo_buf/u_efx_fifo_top/raddr[10] , 
        \u_afifo_buf/u_efx_fifo_top/raddr[11] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] , 
        n769, n770, n771, n772, n773, n774, n775, n776, n777, 
        n778, n779, n780, n781, n782, n783, n784, n785, n786, 
        n787, n788, n789, n790, n791, n792, n793, n794, n795, 
        n796, n797, n798, n799, n800, n801, n802, n803, \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13] , 
        n900, n901, \u_scaler_gray/vs_cnt[0] , n904, n905, tvsync_o, 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] , \u_scaler_gray/tvalid_o_r , 
        n911, n912, \u_scaler_gray/u0_data_stream_ctr/w_addra[0] , n916, 
        n917, \u_scaler_gray/u0_data_stream_ctr/scaler_st[0] , n919, n920, 
        n921, n922, n923, n924, n925, n926, n927, \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0] , 
        \u_scaler_gray/destx[0] , n930, n931, n932, n933, n934, 
        n935, n936, n937, \u_scaler_gray/desty[0] , n940, n941, 
        n942, n943, n944, n945, n946, n947, n948, n949, n950, 
        n951, n952, n953, n954, n955, n956, n957, n958, n959, 
        n960, n961, n962, \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0] , n965, \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0] , 
        \u_scaler_gray/tdata00[1] , \u_scaler_gray/tdata00[0] , \u_scaler_gray/tdata01[1] , 
        \u_scaler_gray/tdata01[0] , \u_scaler_gray/tdata10[0] , \u_scaler_gray/tdata11[0] , 
        n973, n974, \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] , \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] , n1008, n1009, 
        n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
        n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, 
        n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
        n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, 
        n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[11] , \u_scaler_gray/u0_data_stream_ctr/w_addra[12] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[13] , \u_scaler_gray/u0_data_stream_ctr/w_addra[14] , 
        \u_scaler_gray/u0_data_stream_ctr/w_addra[15] , n1065, n1066, 
        n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
        n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
        n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, 
        n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, 
        n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
        n1107, n1108, n1109, n1110, n1111, \u_scaler_gray/u0_data_stream_ctr/scaler_st[1] , 
        \u_scaler_gray/u0_data_stream_ctr/scaler_st[2] , n1114, n1115, 
        \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1] , \u_scaler_gray/destx[1] , 
        \u_scaler_gray/destx[2] , \u_scaler_gray/destx[3] , \u_scaler_gray/destx[4] , 
        \u_scaler_gray/destx[5] , \u_scaler_gray/destx[6] , \u_scaler_gray/destx[7] , 
        \u_scaler_gray/destx[8] , \u_scaler_gray/destx[9] , \u_scaler_gray/destx[10] , 
        \u_scaler_gray/destx[11] , \u_scaler_gray/destx[12] , \u_scaler_gray/destx[13] , 
        \u_scaler_gray/destx[14] , \u_scaler_gray/destx[15] , n1132, n1133, 
        n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, 
        n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
        n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, 
        n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, 
        n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
        n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, 
        n1182, n1183, \u_scaler_gray/desty[1] , \u_scaler_gray/desty[2] , 
        \u_scaler_gray/desty[3] , \u_scaler_gray/desty[4] , \u_scaler_gray/desty[5] , 
        \u_scaler_gray/desty[6] , \u_scaler_gray/desty[7] , \u_scaler_gray/desty[8] , 
        \u_scaler_gray/desty[9] , \u_scaler_gray/desty[10] , \u_scaler_gray/desty[11] , 
        \u_scaler_gray/desty[12] , \u_scaler_gray/desty[13] , \u_scaler_gray/desty[14] , 
        \u_scaler_gray/desty[15] , n1199, n1200, n1201, n1202, n1203, 
        n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, 
        n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
        n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
        n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
        n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, 
        n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, 
        n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
        n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8] , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10] , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11] , 
        n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
        n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, 
        n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, 
        n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, 
        n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, 
        n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
        n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, 
        n1328, \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1] , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3] , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5] , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7] , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9] , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10] , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11] , 
        n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
        n1359, n1360, \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9] , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11] , \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1] , 
        \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2] , \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] , 
        \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4] , \u_scaler_gray/tvalid , 
        \u_scaler_gray/tdata00[2] , \u_scaler_gray/tdata00[3] , \u_scaler_gray/tdata00[4] , 
        \u_scaler_gray/tdata00[5] , \u_scaler_gray/tdata00[6] , \u_scaler_gray/tdata00[7] , 
        \u_scaler_gray/tdata01[2] , \u_scaler_gray/tdata01[3] , \u_scaler_gray/tdata01[4] , 
        \u_scaler_gray/tdata01[5] , \u_scaler_gray/tdata01[6] , \u_scaler_gray/tdata01[7] , 
        \u_scaler_gray/tdata10[1] , \u_scaler_gray/tdata10[2] , \u_scaler_gray/tdata10[3] , 
        \u_scaler_gray/tdata10[4] , \u_scaler_gray/tdata10[5] , \u_scaler_gray/tdata10[6] , 
        \u_scaler_gray/tdata10[7] , \u_scaler_gray/tdata11[1] , \u_scaler_gray/tdata11[2] , 
        \u_scaler_gray/tdata11[3] , \u_scaler_gray/tdata11[4] , \u_scaler_gray/tdata11[5] , 
        \u_scaler_gray/tdata11[6] , \u_scaler_gray/tdata11[7] , n1396, 
        n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, 
        n1405, n1406, \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13] , 
        \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14] , \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15] , 
        n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, 
        n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, 
        n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
        n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, 
        n1481, n1495, n1496, n1497, n1498, n1499, n1500, n1501, 
        n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
        n1510, n1511, n1512, n1513, n1514, n1515, n1516, \u_scaler_gray/vs_cnt[1] , 
        \u_scaler_gray/vs_cnt[2] , \u_scaler_gray/vs_cnt[3] , \u_scaler_gray/vs_cnt[4] , 
        \u_scaler_gray/vs_cnt[5] , \u_scaler_gray/vs_cnt[6] , \u_scaler_gray/vs_cnt[7] , 
        \u_scaler_gray/vs_cnt[8] , \u_scaler_gray/vs_cnt[9] , \u_scaler_gray/vs_cnt[10] , 
        \u_scaler_gray/vs_cnt[11] , \u_scaler_gray/vs_cnt[12] , \u_scaler_gray/vs_cnt[13] , 
        \u_scaler_gray/vs_cnt[14] , \u_scaler_gray/vs_cnt[15] , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[0] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0] , 
        n1534, n1535, n1536, n1537, \u_scaler_gray/u1_bilinear_gray/srcy_fix[0] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[1] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[2] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[3] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[4] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[5] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[6] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[7] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[8] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[9] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[10] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[11] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[12] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[13] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[14] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[15] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[16] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[17] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[18] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[19] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[20] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[21] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[22] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[23] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[24] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[25] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[26] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[27] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27] , 
        \u_scaler_gray/u1_bilinear_gray/srcx_fix[9] , \u_scaler_gray/u1_bilinear_gray/srcx_fix[10] , 
        \u_scaler_gray/u1_bilinear_gray/srcx_fix[11] , \u_scaler_gray/srcx_int[0] , 
        \u_scaler_gray/srcx_int[1] , \u_scaler_gray/srcx_int[2] , \u_scaler_gray/srcx_int[3] , 
        \u_scaler_gray/srcx_int[4] , \u_scaler_gray/srcx_int[5] , \u_scaler_gray/srcx_int[6] , 
        \u_scaler_gray/srcx_int[7] , \u_scaler_gray/srcx_int[8] , \u_scaler_gray/srcx_int[9] , 
        \u_scaler_gray/srcx_int[10] , \u_scaler_gray/srcx_int[11] , \u_scaler_gray/srcx_int[12] , 
        \u_scaler_gray/srcx_int[13] , \u_scaler_gray/srcx_int[14] , \u_scaler_gray/srcx_int[15] , 
        n1640, n1641, n1642, n1643, \u_scaler_gray/u1_bilinear_gray/srcy_fix[1] , 
        \u_scaler_gray/u1_bilinear_gray/srcy_fix[2] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[3] , 
        \u_scaler_gray/u1_bilinear_gray/srcy_fix[4] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[5] , 
        \u_scaler_gray/u1_bilinear_gray/srcy_fix[6] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[7] , 
        \u_scaler_gray/u1_bilinear_gray/srcy_fix[8] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[9] , 
        \u_scaler_gray/u1_bilinear_gray/srcy_fix[10] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[11] , 
        \u_scaler_gray/srcy_int[0] , \u_scaler_gray/srcy_int[1] , \u_scaler_gray/srcy_int[2] , 
        \u_scaler_gray/srcy_int[3] , \u_scaler_gray/srcy_int[4] , \u_scaler_gray/srcy_int[5] , 
        \u_scaler_gray/srcy_int[6] , \u_scaler_gray/srcy_int[7] , \u_scaler_gray/srcy_int[8] , 
        \u_scaler_gray/srcy_int[9] , \u_scaler_gray/srcy_int[10] , \u_scaler_gray/srcy_int[11] , 
        \u_scaler_gray/srcy_int[12] , \u_scaler_gray/srcy_int[13] , \u_scaler_gray/srcy_int[14] , 
        \u_scaler_gray/srcy_int[15] , n1671, n1672, n1673, n1674, 
        n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
        n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, 
        n1691, n1692, n1693, \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0] , 
        n1713, n1714, n1719, n1720, n1721, n1722, n1723, n1724, 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11] , 
        n1739, n1740, n1769, n1770, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[11] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[12] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[13] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[14] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[15] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[16] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[17] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[18] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[19] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[20] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[21] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[22] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[23] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[11] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[12] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[13] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[14] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[15] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[16] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[17] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[18] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[19] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[20] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[21] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[22] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[23] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[11] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[12] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[13] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[14] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[15] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[16] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[17] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[18] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[19] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[20] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[21] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[22] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[23] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[11] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[12] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[13] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[14] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[15] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[16] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[17] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[18] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[19] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[20] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[21] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[22] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[23] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10] , 
        \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[5] , 
        n1908, n1909, n1910, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[4] , 
        n1913, n1914, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[3] , 
        \tdata_o[0] , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[0] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9] , 
        \tdata_o[1] , \tdata_o[2] , \tdata_o[3] , \tdata_o[4] , \tdata_o[5] , 
        \tdata_o[6] , \tdata_o[7] , n2054, n2055, n2056, n2057, 
        n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, 
        n2066, n2067, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[1] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[2] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[3] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[4] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[5] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[6] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[7] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[8] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[9] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[10] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[11] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[12] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[13] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[14] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[15] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[16] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[17] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[18] , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[19] , 
        n2107, n2108, n2109, n2110, \u_axi4_ctrl/wframe_vsync_dly[0] , 
        n2112, n2113, \u_axi4_ctrl/wframe_index[1] , n2115, n2116, 
        \u_axi4_ctrl/rframe_vsync_dly[0] , n2119, n2120, \u_axi4_ctrl/wframe_index[0] , 
        n2122, n2123, n2124, n2125, n2126, n2127, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , 
        \u_axi4_ctrl/rframe_index[0] , n2132, n2133, n2134, \u_axi4_ctrl/state[0] , 
        n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, 
        n2144, n2145, \u_axi4_ctrl/wframe_vsync_dly[1] , n2147, n2148, 
        n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, 
        n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, 
        n2166, n2167, \u_axi4_ctrl/wframe_vsync_dly[3] , n2169, n2170, 
        n2187, n2188, n2189, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , n2224, n2225, 
        n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, 
        n2234, n2235, n2269, n2270, n2271, n2272, n2291, n2292, 
        n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, 
        n2304, n2305, \u_axi4_ctrl/wdata_cnt_dly[0] , \u_axi4_ctrl/rdata_cnt_dly[1] , 
        \u_axi4_ctrl/rdata_cnt_dly[0] , \u_axi4_ctrl/rframe_vsync_dly[3] , 
        n2312, n2313, n2314, n2315, n2316, \u_axi4_ctrl/rfifo_wenb , 
        n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, 
        n2328, n2329, n2330, n2331, \u_axi4_ctrl/rfifo_wdata[0] , 
        n2334, n2335, n2336, n2337, n2338, n2339, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/wfifo_empty , 
        n2343, n2344, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
        n2346, n2347, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] , 
        n2349, n2350, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] , 
        n2352, n2353, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , 
        n2355, n2356, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , 
        n2367, n2369, n2370, n2371, n2372, n2373, n2374, n2375, 
        n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] , 
        n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, 
        n2400, n2401, n2402, n2403, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] , 
        n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
        n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, 
        n2499, n2510, n2511, n2512, n2513, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] , 
        \u_axi4_ctrl/rfifo_empty , n2517, n2518, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] , 
        n2520, n2521, n2522, n2523, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] , 
        n2527, n2528, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] , 
        n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
        n2545, n2546, n2547, n2548, n2549, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] , 
        n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, 
        n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, 
        n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, 
        n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, 
        n2594, n2595, n2596, n2597, n2598, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] , 
        n2679, n2680, n2681, n2682, n2683, n2684, \u_axi4_ctrl/rframe_index[1] , 
        n2686, n2687, \u_axi4_ctrl/state[1] , \u_axi4_ctrl/state[2] , 
        n2690, n2691, n2692, n2693, \u_axi4_ctrl/awaddr[10] , \u_axi4_ctrl/awaddr[11] , 
        \u_axi4_ctrl/awaddr[12] , \u_axi4_ctrl/awaddr[13] , \u_axi4_ctrl/awaddr[14] , 
        \u_axi4_ctrl/awaddr[15] , \u_axi4_ctrl/awaddr[16] , \u_axi4_ctrl/awaddr[17] , 
        \u_axi4_ctrl/awaddr[18] , \u_axi4_ctrl/awaddr[19] , \u_axi4_ctrl/awaddr[20] , 
        \u_axi4_ctrl/awaddr[21] , \u_axi4_ctrl/awaddr[22] , \u_axi4_ctrl/awaddr[23] , 
        n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, 
        n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, 
        n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, 
        n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, 
        n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, 
        n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, 
        n2776, n2777, \u_axi4_ctrl/araddr[10] , \u_axi4_ctrl/araddr[11] , 
        \u_axi4_ctrl/araddr[12] , \u_axi4_ctrl/araddr[13] , \u_axi4_ctrl/araddr[14] , 
        \u_axi4_ctrl/araddr[15] , \u_axi4_ctrl/araddr[16] , \u_axi4_ctrl/araddr[17] , 
        \u_axi4_ctrl/araddr[18] , \u_axi4_ctrl/araddr[19] , \u_axi4_ctrl/araddr[20] , 
        \u_axi4_ctrl/araddr[21] , \u_axi4_ctrl/araddr[22] , \u_axi4_ctrl/araddr[23] , 
        n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, 
        n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, 
        n2808, n2809, n2810, n2811, n2812, n2855, n2856, n2857, 
        n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, 
        n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
        n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, 
        n2882, \u_axi4_ctrl/wdata_cnt_dly[1] , \u_axi4_ctrl/wdata_cnt_dly[2] , 
        \u_axi4_ctrl/wdata_cnt_dly[3] , \u_axi4_ctrl/wdata_cnt_dly[4] , 
        \u_axi4_ctrl/wdata_cnt_dly[5] , \u_axi4_ctrl/wdata_cnt_dly[6] , 
        \u_axi4_ctrl/wdata_cnt_dly[7] , \u_axi4_ctrl/wdata_cnt_dly[8] , 
        \u_axi4_ctrl/rdata_cnt_dly[2] , \u_axi4_ctrl/rdata_cnt_dly[3] , 
        \u_axi4_ctrl/rdata_cnt_dly[4] , \u_axi4_ctrl/rdata_cnt_dly[5] , 
        \u_axi4_ctrl/rdata_cnt_dly[6] , \u_axi4_ctrl/rdata_cnt_dly[7] , 
        \u_axi4_ctrl/rdata_cnt_dly[8] , n2898, n2899, n2900, n2901, 
        \u_axi4_ctrl/rfifo_wdata[1] , \u_axi4_ctrl/rfifo_wdata[2] , \u_axi4_ctrl/rfifo_wdata[3] , 
        \u_axi4_ctrl/rfifo_wdata[4] , \u_axi4_ctrl/rfifo_wdata[5] , \u_axi4_ctrl/rfifo_wdata[6] , 
        \u_axi4_ctrl/rfifo_wdata[7] , \u_axi4_ctrl/rfifo_wdata[8] , \u_axi4_ctrl/rfifo_wdata[9] , 
        \u_axi4_ctrl/rfifo_wdata[10] , \u_axi4_ctrl/rfifo_wdata[11] , \u_axi4_ctrl/rfifo_wdata[12] , 
        \u_axi4_ctrl/rfifo_wdata[13] , \u_axi4_ctrl/rfifo_wdata[14] , \u_axi4_ctrl/rfifo_wdata[15] , 
        \u_axi4_ctrl/rfifo_wdata[16] , \u_axi4_ctrl/rfifo_wdata[17] , \u_axi4_ctrl/rfifo_wdata[18] , 
        \u_axi4_ctrl/rfifo_wdata[19] , \u_axi4_ctrl/rfifo_wdata[20] , \u_axi4_ctrl/rfifo_wdata[21] , 
        \u_axi4_ctrl/rfifo_wdata[22] , \u_axi4_ctrl/rfifo_wdata[23] , \u_axi4_ctrl/rfifo_wdata[24] , 
        \u_axi4_ctrl/rfifo_wdata[25] , \u_axi4_ctrl/rfifo_wdata[26] , \u_axi4_ctrl/rfifo_wdata[27] , 
        \u_axi4_ctrl/rfifo_wdata[28] , \u_axi4_ctrl/rfifo_wdata[29] , \u_axi4_ctrl/rfifo_wdata[30] , 
        \u_axi4_ctrl/rfifo_wdata[31] , \u_axi4_ctrl/rfifo_wdata[32] , \u_axi4_ctrl/rfifo_wdata[33] , 
        \u_axi4_ctrl/rfifo_wdata[34] , \u_axi4_ctrl/rfifo_wdata[35] , \u_axi4_ctrl/rfifo_wdata[36] , 
        \u_axi4_ctrl/rfifo_wdata[37] , \u_axi4_ctrl/rfifo_wdata[38] , \u_axi4_ctrl/rfifo_wdata[39] , 
        \u_axi4_ctrl/rfifo_wdata[40] , \u_axi4_ctrl/rfifo_wdata[41] , \u_axi4_ctrl/rfifo_wdata[42] , 
        \u_axi4_ctrl/rfifo_wdata[43] , \u_axi4_ctrl/rfifo_wdata[44] , \u_axi4_ctrl/rfifo_wdata[45] , 
        \u_axi4_ctrl/rfifo_wdata[46] , \u_axi4_ctrl/rfifo_wdata[47] , \u_axi4_ctrl/rfifo_wdata[48] , 
        \u_axi4_ctrl/rfifo_wdata[49] , \u_axi4_ctrl/rfifo_wdata[50] , \u_axi4_ctrl/rfifo_wdata[51] , 
        \u_axi4_ctrl/rfifo_wdata[52] , \u_axi4_ctrl/rfifo_wdata[53] , \u_axi4_ctrl/rfifo_wdata[54] , 
        \u_axi4_ctrl/rfifo_wdata[55] , \u_axi4_ctrl/rfifo_wdata[56] , \u_axi4_ctrl/rfifo_wdata[57] , 
        \u_axi4_ctrl/rfifo_wdata[58] , \u_axi4_ctrl/rfifo_wdata[59] , \u_axi4_ctrl/rfifo_wdata[60] , 
        \u_axi4_ctrl/rfifo_wdata[61] , \u_axi4_ctrl/rfifo_wdata[62] , \u_axi4_ctrl/rfifo_wdata[63] , 
        \u_axi4_ctrl/rfifo_wdata[64] , \u_axi4_ctrl/rfifo_wdata[65] , \u_axi4_ctrl/rfifo_wdata[66] , 
        \u_axi4_ctrl/rfifo_wdata[67] , \u_axi4_ctrl/rfifo_wdata[68] , \u_axi4_ctrl/rfifo_wdata[69] , 
        \u_axi4_ctrl/rfifo_wdata[70] , \u_axi4_ctrl/rfifo_wdata[71] , \u_axi4_ctrl/rfifo_wdata[72] , 
        \u_axi4_ctrl/rfifo_wdata[73] , \u_axi4_ctrl/rfifo_wdata[74] , \u_axi4_ctrl/rfifo_wdata[75] , 
        \u_axi4_ctrl/rfifo_wdata[76] , \u_axi4_ctrl/rfifo_wdata[77] , \u_axi4_ctrl/rfifo_wdata[78] , 
        \u_axi4_ctrl/rfifo_wdata[79] , \u_axi4_ctrl/rfifo_wdata[80] , \u_axi4_ctrl/rfifo_wdata[81] , 
        \u_axi4_ctrl/rfifo_wdata[82] , \u_axi4_ctrl/rfifo_wdata[83] , \u_axi4_ctrl/rfifo_wdata[84] , 
        \u_axi4_ctrl/rfifo_wdata[85] , \u_axi4_ctrl/rfifo_wdata[86] , \u_axi4_ctrl/rfifo_wdata[87] , 
        \u_axi4_ctrl/rfifo_wdata[88] , \u_axi4_ctrl/rfifo_wdata[89] , \u_axi4_ctrl/rfifo_wdata[90] , 
        \u_axi4_ctrl/rfifo_wdata[91] , \u_axi4_ctrl/rfifo_wdata[92] , \u_axi4_ctrl/rfifo_wdata[93] , 
        \u_axi4_ctrl/rfifo_wdata[94] , \u_axi4_ctrl/rfifo_wdata[95] , \u_axi4_ctrl/rfifo_wdata[96] , 
        \u_axi4_ctrl/rfifo_wdata[97] , \u_axi4_ctrl/rfifo_wdata[98] , \u_axi4_ctrl/rfifo_wdata[99] , 
        \u_axi4_ctrl/rfifo_wdata[100] , \u_axi4_ctrl/rfifo_wdata[101] , 
        \u_axi4_ctrl/rfifo_wdata[102] , \u_axi4_ctrl/rfifo_wdata[103] , 
        \u_axi4_ctrl/rfifo_wdata[104] , \u_axi4_ctrl/rfifo_wdata[105] , 
        \u_axi4_ctrl/rfifo_wdata[106] , \u_axi4_ctrl/rfifo_wdata[107] , 
        \u_axi4_ctrl/rfifo_wdata[108] , \u_axi4_ctrl/rfifo_wdata[109] , 
        \u_axi4_ctrl/rfifo_wdata[110] , \u_axi4_ctrl/rfifo_wdata[111] , 
        \u_axi4_ctrl/rfifo_wdata[112] , \u_axi4_ctrl/rfifo_wdata[113] , 
        \u_axi4_ctrl/rfifo_wdata[114] , \u_axi4_ctrl/rfifo_wdata[115] , 
        \u_axi4_ctrl/rfifo_wdata[116] , \u_axi4_ctrl/rfifo_wdata[117] , 
        \u_axi4_ctrl/rfifo_wdata[118] , \u_axi4_ctrl/rfifo_wdata[119] , 
        \u_axi4_ctrl/rfifo_wdata[120] , \u_axi4_ctrl/rfifo_wdata[121] , 
        \u_axi4_ctrl/rfifo_wdata[122] , \u_axi4_ctrl/rfifo_wdata[123] , 
        \u_axi4_ctrl/rfifo_wdata[124] , \u_axi4_ctrl/rfifo_wdata[125] , 
        \u_axi4_ctrl/rfifo_wdata[126] , \u_axi4_ctrl/rfifo_wdata[127] , 
        n3029, n3030, n3031, n3032, \u_lcd_driver/vcnt[0] , lcd_hs, 
        n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, 
        lcd_de, n3045, n3046, n3047, n3048, \u_lcd_driver/r_lcd_dv , 
        \u_lcd_driver/hcnt[0] , n3052, n3053, n3054, n3055, \u_lcd_driver/vcnt[1] , 
        \u_lcd_driver/vcnt[2] , \u_lcd_driver/vcnt[3] , \u_lcd_driver/vcnt[4] , 
        \u_lcd_driver/vcnt[5] , \u_lcd_driver/vcnt[6] , \u_lcd_driver/vcnt[7] , 
        \u_lcd_driver/vcnt[8] , \u_lcd_driver/vcnt[9] , \u_lcd_driver/vcnt[10] , 
        \u_lcd_driver/vcnt[11] , n3067, n3068, n3069, n3070, n3071, 
        n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, 
        n3080, n3081, n3082, \u_lcd_driver/r_lcd_rgb[5] , \u_lcd_driver/hcnt[1] , 
        \u_lcd_driver/hcnt[2] , \u_lcd_driver/hcnt[3] , \u_lcd_driver/hcnt[4] , 
        \u_lcd_driver/hcnt[5] , \u_lcd_driver/hcnt[6] , \u_lcd_driver/hcnt[7] , 
        \u_lcd_driver/hcnt[8] , \u_lcd_driver/hcnt[9] , \u_lcd_driver/hcnt[10] , 
        \u_lcd_driver/hcnt[11] , n3195, n3196, \w_hdmi_txd0[0] , \u_rgb2dvi/enc_0/acc[0] , 
        n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, 
        n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, 
        n3223, n3224, n3225, n3226, n3227, \w_hdmi_txd0[1] , \w_hdmi_txd0[2] , 
        \w_hdmi_txd0[3] , \w_hdmi_txd0[4] , \w_hdmi_txd0[5] , \w_hdmi_txd0[6] , 
        \w_hdmi_txd0[7] , \w_hdmi_txd0[8] , \w_hdmi_txd0[9] , \u_rgb2dvi/enc_0/acc[1] , 
        \u_rgb2dvi/enc_0/acc[2] , \u_rgb2dvi/enc_0/acc[3] , \u_rgb2dvi/enc_0/acc[4] , 
        n3254, n3255, \w_hdmi_txd1[0] , \u_rgb2dvi/enc_1/acc[0] , n3284, 
        n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, 
        n3293, n3294, n3295, n3296, n3297, n3298, n3299, \w_hdmi_txd1[1] , 
        \w_hdmi_txd1[2] , \w_hdmi_txd1[3] , \w_hdmi_txd1[4] , \w_hdmi_txd1[5] , 
        \w_hdmi_txd1[6] , \w_hdmi_txd1[7] , \w_hdmi_txd1[8] , \w_hdmi_txd1[9] , 
        n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, 
        \u_rgb2dvi/enc_1/acc[1] , \u_rgb2dvi/enc_1/acc[2] , \u_rgb2dvi/enc_1/acc[3] , 
        \u_rgb2dvi/enc_1/acc[4] , n3321, n3322, n3323, n3324, n3325, 
        n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, 
        n3334, n3335, n3336, \w_hdmi_txd2[0] , n3338, n3339, \u_rgb2dvi/enc_2/acc[0] , 
        n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, 
        n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
        n3357, n3358, n3359, n3360, n3361, \w_hdmi_txd2[1] , \w_hdmi_txd2[2] , 
        \w_hdmi_txd2[3] , \w_hdmi_txd2[4] , \w_hdmi_txd2[5] , \w_hdmi_txd2[6] , 
        \w_hdmi_txd2[7] , \w_hdmi_txd2[9] , n3370, n3371, n3372, n3373, 
        n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, 
        n3382, n3383, \u_rgb2dvi/enc_2/acc[1] , \u_rgb2dvi/enc_2/acc[2] , 
        \u_rgb2dvi/enc_2/acc[3] , \u_rgb2dvi/enc_2/acc[4] , n3388, n3389, 
        n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, 
        n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, 
        n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, 
        n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, 
        n3422, n3423, n3424, n3426, n3427, n3428, n3429, n3430, 
        \r_hdmi_tx0_o[5] , \r_hdmi_tx0_o[6] , \r_hdmi_tx0_o[7] , \r_hdmi_tx0_o[8] , 
        \r_hdmi_tx0_o[9] , \r_hdmi_tx1_o[5] , \r_hdmi_tx1_o[6] , \r_hdmi_tx1_o[7] , 
        \r_hdmi_tx1_o[8] , \r_hdmi_tx1_o[9] , \r_hdmi_tx2_o[5] , \r_hdmi_tx2_o[6] , 
        \r_hdmi_tx2_o[7] , \r_hdmi_tx2_o[9] , \PowerOnResetCnt[1] , \PowerOnResetCnt[2] , 
        \PowerOnResetCnt[3] , \PowerOnResetCnt[4] , \PowerOnResetCnt[5] , 
        \PowerOnResetCnt[6] , \PowerOnResetCnt[7] , n3465, n3466, n3467, 
        n3468, n3469, n3470, n3471, n3472, n3473, n3474, \reduce_nand_9/n7 , 
        DdrInitDone, \Axi0ResetReg[2] , \cmos_frame_Gray[2] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n15 , \U0_DDR_Reset/u_ddr_reset_sequencer/equal_21/n3 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] , \U0_DDR_Reset/u_ddr_reset_sequencer/n92 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] , \U0_DDR_Reset/u_ddr_reset_sequencer/n91 , 
        \u_i2c_timing_ctrl_16reg_16bit/n137 , \u_i2c_timing_ctrl_16reg_16bit/next_state[1] , 
        \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en , \u_i2c_timing_ctrl_16reg_16bit/next_state[0] , 
        \u_i2c_timing_ctrl_16reg_16bit/n138 , \u_i2c_timing_ctrl_16reg_16bit/n139 , 
        \u_i2c_timing_ctrl_16reg_16bit/n140 , \u_i2c_timing_ctrl_16reg_16bit/n205 , 
        \u_i2c_timing_ctrl_16reg_16bit/n846 , \u_i2c_timing_ctrl_16reg_16bit/n122 , 
        \u_i2c_timing_ctrl_16reg_16bit/n123 , \u_i2c_timing_ctrl_16reg_16bit/n124 , 
        \u_i2c_timing_ctrl_16reg_16bit/n125 , \u_i2c_timing_ctrl_16reg_16bit/n126 , 
        \u_i2c_timing_ctrl_16reg_16bit/n127 , \u_i2c_timing_ctrl_16reg_16bit/n128 , 
        \u_i2c_timing_ctrl_16reg_16bit/n129 , \u_i2c_timing_ctrl_16reg_16bit/n130 , 
        \u_i2c_timing_ctrl_16reg_16bit/n131 , \u_i2c_timing_ctrl_16reg_16bit/n132 , 
        \u_i2c_timing_ctrl_16reg_16bit/n133 , \u_i2c_timing_ctrl_16reg_16bit/n134 , 
        \u_i2c_timing_ctrl_16reg_16bit/n135 , \u_i2c_timing_ctrl_16reg_16bit/n136 , 
        \u_i2c_timing_ctrl_16reg_16bit/n500 , ceg_net552, \u_i2c_timing_ctrl_16reg_16bit/n509 , 
        ceg_net664, \u_i2c_timing_ctrl_16reg_16bit/n567 , \u_i2c_timing_ctrl_16reg_16bit/n570 , 
        \u_i2c_timing_ctrl_16reg_16bit/n573 , \u_i2c_timing_ctrl_16reg_16bit/n576 , 
        \u_i2c_timing_ctrl_16reg_16bit/n579 , \u_i2c_timing_ctrl_16reg_16bit/n581 , 
        \u_i2c_timing_ctrl_16reg_16bit/n7 , \u_i2c_timing_ctrl_16reg_16bit/n495 , 
        ceg_net632, \u_i2c_timing_ctrl_16reg_16bit/next_state[2] , \u_i2c_timing_ctrl_16reg_16bit/next_state[3] , 
        \u_i2c_timing_ctrl_16reg_16bit/next_state[4] , \u_i2c_timing_ctrl_16reg_16bit/n204 , 
        \u_i2c_timing_ctrl_16reg_16bit/n203 , \u_i2c_timing_ctrl_16reg_16bit/n202 , 
        \u_i2c_timing_ctrl_16reg_16bit/n201 , \u_i2c_timing_ctrl_16reg_16bit/n200 , 
        \u_i2c_timing_ctrl_16reg_16bit/n199 , \u_i2c_timing_ctrl_16reg_16bit/n198 , 
        \u_i2c_timing_ctrl_16reg_16bit/n499 , \u_i2c_timing_ctrl_16reg_16bit/n498 , 
        \u_i2c_timing_ctrl_16reg_16bit/n497 , \u_i2c_timing_ctrl_16reg_16bit/n508 , 
        \u_i2c_timing_ctrl_16reg_16bit/n507 , \u_i2c_timing_ctrl_16reg_16bit/n506 , 
        \u_i2c_timing_ctrl_16reg_16bit/n505 , \u_i2c_timing_ctrl_16reg_16bit/n504 , 
        \u_i2c_timing_ctrl_16reg_16bit/n503 , \u_i2c_timing_ctrl_16reg_16bit/n502 , 
        n3881, n3884, n3887, n3890, n3895, n3898, n3901, n3904, 
        n3913, n3916, n3919, n3920, n3923, n3926, n3932, n3935, 
        n3938, n3941, \u_CMOS_Capture_RAW_Gray/n127 , ceg_net152, \u_CMOS_Capture_RAW_Gray/n160 , 
        ceg_net158, \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7] , \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6] , 
        \u_CMOS_Capture_RAW_Gray/n171 , \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1] , 
        \u_CMOS_Capture_RAW_Gray/n126 , \u_CMOS_Capture_RAW_Gray/n125 , 
        \u_CMOS_Capture_RAW_Gray/n124 , \u_CMOS_Capture_RAW_Gray/n123 , 
        \u_CMOS_Capture_RAW_Gray/n122 , \u_CMOS_Capture_RAW_Gray/n121 , 
        \u_CMOS_Capture_RAW_Gray/n120 , \u_CMOS_Capture_RAW_Gray/n119 , 
        \u_CMOS_Capture_RAW_Gray/n118 , \u_CMOS_Capture_RAW_Gray/n117 , 
        \u_CMOS_Capture_RAW_Gray/n116 , \u_CMOS_Capture_RAW_Gray/n159 , 
        n4132, n4135, n4138, cmos_frame_href, \u_sensor_frame_count/n66 , 
        \u_sensor_frame_count/n67 , \u_sensor_frame_count/n68 , \u_sensor_frame_count/n69 , 
        n4176, \u_sensor_frame_count/n70 , \u_sensor_frame_count/n71 , 
        \u_sensor_frame_count/n74 , \u_sensor_frame_count/cmos_fps_cnt[1] , 
        \u_sensor_frame_count/n141 , ceg_net200, \u_sensor_frame_count/n72 , 
        \u_sensor_frame_count/n73 , \u_sensor_frame_count/n75 , \cmos_frame_Gray[0] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 , \u_sensor_frame_count/n110 , 
        \u_sensor_frame_count/n65 , \u_sensor_frame_count/n64 , \u_sensor_frame_count/n63 , 
        \u_sensor_frame_count/n62 , \u_sensor_frame_count/n61 , \u_sensor_frame_count/n60 , 
        \u_sensor_frame_count/n59 , \u_sensor_frame_count/n58 , \u_sensor_frame_count/n57 , 
        \u_sensor_frame_count/n56 , \u_sensor_frame_count/n55 , \u_sensor_frame_count/n54 , 
        \u_sensor_frame_count/n53 , \u_sensor_frame_count/n52 , \u_sensor_frame_count/n51 , 
        \u_sensor_frame_count/n50 , \u_sensor_frame_count/n49 , \u_sensor_frame_count/n48 , 
        n4211, \u_sensor_frame_count/n140 , \u_sensor_frame_count/n139 , 
        \u_sensor_frame_count/n138 , \u_sensor_frame_count/n137 , \u_sensor_frame_count/n136 , 
        \u_sensor_frame_count/n135 , \u_sensor_frame_count/n134 , \u_sensor_frame_count/n133 , 
        n4222, n4225, \u_afifo_buf/u_efx_fifo_top/raddr[12] , \u_afifo_buf/u_efx_fifo_top/rd_en_int , 
        \cmos_frame_Gray[1] , \cmos_frame_Gray[3] , \cmos_frame_Gray[4] , 
        \cmos_frame_Gray[5] , \cmos_frame_Gray[6] , \cmos_frame_Gray[7] , 
        \u_afifo_buf/u_efx_fifo_top/wr_en_int , ceg_net219, n4296, \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[13] , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[12] , 
        ceg_net226, \u_scaler_gray/n150 , ceg_net229, \u_scaler_gray/u0_data_stream_ctr/w_image_tlast , 
        \u_scaler_gray/u0_data_stream_ctr/n1703 , tvalid_o, \u_scaler_gray/u0_data_stream_ctr/n1704 , 
        \u_scaler_gray/u0_data_stream_ctr/n432 , \u_scaler_gray/u0_data_stream_ctr/n2156 , 
        ceg_net526, \u_scaler_gray/u0_data_stream_ctr/equal_59/n5 , \u_scaler_gray/u0_data_stream_ctr/n1712 , 
        \u_scaler_gray/u0_data_stream_ctr/r_image_tlast , \u_scaler_gray/u0_data_stream_ctr/n1713 , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
        \tdata_i[6] , \u_scaler_gray/u0_data_stream_ctr/n903 , \tdata_i[1] , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
        \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
        \u_scaler_gray/u0_data_stream_ctr/n1702 , \u_scaler_gray/u0_data_stream_ctr/n431 , 
        \u_scaler_gray/u0_data_stream_ctr/n430 , \u_scaler_gray/u0_data_stream_ctr/n2073 , 
        \u_scaler_gray/u0_data_stream_ctr/n1161 , \u_scaler_gray/u0_data_stream_ctr/n1160 , 
        \u_scaler_gray/u0_data_stream_ctr/n1159 , \u_scaler_gray/u0_data_stream_ctr/n885 , 
        \u_scaler_gray/u0_data_stream_ctr/n884 , \u_scaler_gray/u0_data_stream_ctr/n883 , 
        \u_scaler_gray/u0_data_stream_ctr/n882 , \u_scaler_gray/u0_data_stream_ctr/n881 , 
        \u_scaler_gray/u0_data_stream_ctr/n880 , \u_scaler_gray/u0_data_stream_ctr/n879 , 
        \u_scaler_gray/u0_data_stream_ctr/n1179 , \u_scaler_gray/u0_data_stream_ctr/n1178 , 
        \u_scaler_gray/u0_data_stream_ctr/n1177 , \u_scaler_gray/u0_data_stream_ctr/n1176 , 
        \u_scaler_gray/u0_data_stream_ctr/n1196 , \u_scaler_gray/u0_data_stream_ctr/n1195 , 
        \u_scaler_gray/u0_data_stream_ctr/n1194 , \u_scaler_gray/u0_data_stream_ctr/n1193 , 
        \u_scaler_gray/u0_data_stream_ctr/n1212 , \u_scaler_gray/u0_data_stream_ctr/n1211 , 
        \u_scaler_gray/u0_data_stream_ctr/n1210 , \tdata_i[5] , \tdata_i[7] , 
        \tdata_i[4] , \tdata_i[2] , \tdata_i[3] , \tdata_i[0] , \u_scaler_gray/n129 , 
        \u_scaler_gray/n128 , \u_scaler_gray/n127 , \u_scaler_gray/n126 , 
        \u_scaler_gray/n125 , \u_scaler_gray/n124 , \u_scaler_gray/n123 , 
        \u_scaler_gray/n122 , \u_scaler_gray/n121 , \u_scaler_gray/n120 , 
        \u_scaler_gray/n119 , \u_scaler_gray/n118 , \u_scaler_gray/n117 , 
        \u_scaler_gray/n116 , \u_scaler_gray/n115 , \hdmi_clk1x_i~O , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n462 , \hdmi_clk2x_i~O , 
        \cmos_pclk~O , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10] , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n335 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n334 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n333 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n332 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n331 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n330 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n329 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n328 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n327 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n326 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n325 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n324 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n323 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n322 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n321 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n320 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n319 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n318 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n317 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n461 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n460 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n459 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n458 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n457 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n456 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n455 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n454 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n453 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n452 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n451 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n450 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n449 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n448 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n447 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n446 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n445 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n444 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n443 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n442 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n441 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n440 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n439 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n438 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n437 , 
        \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n436 , \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n435 , 
        n7562, n7563, n7564, n7565, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n344 , 
        n7566, n7567, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 , 
        n7568, n7569, n7570, n7571, n7572, n7574, n7575, n7576, 
        n7577, n7578, n7579, \Axi_Clk~O , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n343 , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n342 , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n341 , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n340 , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n339 , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n338 , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n337 , 
        \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n336 , \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n335 , 
        \u_axi4_ctrl/n316 , \u_axi4_ctrl/equal_38/n3 , lcd_vs, \u_axi4_ctrl/n1469 , 
        \u_axi4_ctrl/n317 , \u_axi4_ctrl/n336 , \u_axi4_ctrl/equal_47/n3 , 
        \u_axi4_ctrl/n389 , \u_axi4_ctrl/n405 , \u_axi4_ctrl/n1476 , \u_axi4_ctrl/wframe_vsync_dly[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int , 
        \u_axi4_ctrl/n363 , \u_axi4_ctrl/n1544 , \u_axi4_ctrl/n379 , \u_axi4_ctrl/rframe_vsync_dly[2] , 
        \u_axi4_ctrl/rframe_vsync_dly[1] , ceg_net289, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] , 
        n5870, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] , 
        ceg_net296, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] , 
        \u_axi4_ctrl/n335 , \u_axi4_ctrl/n1610 , \u_axi4_ctrl/n1617 , 
        \u_axi4_ctrl/n387 , \u_axi4_ctrl/n369 , n6308, n6311, n6314, 
        n6317, n6320, n6323, n6326, n6329, n6332, n6335, n6338, 
        n6341, \u_axi4_ctrl/n381 , \u_axi4_ctrl/n1478 , \u_axi4_ctrl/n697 , 
        ceg_net401, \u_axi4_ctrl/n696 , \u_axi4_ctrl/n695 , \u_axi4_ctrl/n694 , 
        \u_axi4_ctrl/n693 , \u_axi4_ctrl/n692 , \u_axi4_ctrl/n691 , \u_axi4_ctrl/n690 , 
        \u_axi4_ctrl/n689 , \u_axi4_ctrl/n688 , \u_axi4_ctrl/n687 , \u_axi4_ctrl/n686 , 
        \u_axi4_ctrl/n685 , \u_axi4_ctrl/n684 , \u_axi4_ctrl/n683 , \u_axi4_ctrl/n682 , 
        \u_axi4_ctrl/n1499 , \u_axi4_ctrl/n1504 , \u_axi4_ctrl/n1509 , 
        \u_axi4_ctrl/n1514 , \u_axi4_ctrl/n1519 , \u_axi4_ctrl/n1524 , 
        \u_axi4_ctrl/n1529 , \u_axi4_ctrl/n1534 , \u_axi4_ctrl/n1549 , 
        \u_axi4_ctrl/n1554 , \u_axi4_ctrl/n1559 , \u_axi4_ctrl/n1564 , 
        \u_axi4_ctrl/n1569 , \u_axi4_ctrl/n1574 , \u_axi4_ctrl/n1579 , 
        \u_lcd_driver/n83 , \u_lcd_driver/equal_17/n23 , \u_lcd_driver/n35 , 
        \u_lcd_driver/n97 , \u_lcd_driver/n125 , \lcd_data[0] , \u_lcd_driver/n133 , 
        \u_lcd_driver/n34 , \u_lcd_driver/n82 , \u_lcd_driver/n81 , \u_lcd_driver/n80 , 
        \u_lcd_driver/n79 , \u_lcd_driver/n78 , \u_lcd_driver/n77 , \u_lcd_driver/n76 , 
        \u_lcd_driver/n75 , \u_lcd_driver/n74 , \u_lcd_driver/n73 , \u_lcd_driver/n72 , 
        \lcd_data[1] , \lcd_data[2] , \lcd_data[3] , \lcd_data[4] , 
        \lcd_data[5] , \lcd_data[6] , \lcd_data[7] , \u_lcd_driver/n33 , 
        \u_lcd_driver/n32 , \u_lcd_driver/n31 , \u_lcd_driver/n30 , \u_lcd_driver/n29 , 
        \u_lcd_driver/n28 , \u_lcd_driver/n27 , \u_lcd_driver/n26 , \u_lcd_driver/n25 , 
        \u_lcd_driver/n24 , \u_lcd_driver/n23 , \u_rgb2dvi/enc_0/n869 , 
        \u_rgb2dvi/enc_0/n764 , \u_rgb2dvi/enc_0/n770 , \u_rgb2dvi/enc_0/n776 , 
        \u_rgb2dvi/enc_0/n782 , \u_rgb2dvi/enc_0/n788 , \u_rgb2dvi/enc_0/n794 , 
        \u_rgb2dvi/enc_0/n800 , \u_rgb2dvi/enc_0/n806 , \u_rgb2dvi/enc_0/n812 , 
        \u_rgb2dvi/enc_1/q_out[0] , \u_rgb2dvi/enc_1/q_out[1] , \u_rgb2dvi/enc_1/q_out[2] , 
        \u_rgb2dvi/enc_1/q_out[3] , \u_rgb2dvi/enc_1/q_out[4] , \u_rgb2dvi/enc_1/q_out[5] , 
        \u_rgb2dvi/enc_1/q_out[6] , \u_rgb2dvi/enc_1/q_out[7] , \u_rgb2dvi/enc_0/n103 , 
        \u_rgb2dvi/enc_1/q_out[9] , n6895, \u_rgb2dvi/enc_2/q_out[0] , 
        \u_rgb2dvi/enc_2/q_out[1] , \u_rgb2dvi/enc_2/q_out[2] , \u_rgb2dvi/enc_2/q_out[3] , 
        \u_rgb2dvi/enc_2/q_out[4] , \u_rgb2dvi/enc_2/q_out[5] , \u_rgb2dvi/enc_2/q_out[6] , 
        \u_rgb2dvi/enc_2/q_out[7] , \u_rgb2dvi/enc_2/q_out[9] , \r_hdmi_txc_o[9] , 
        n591, n590, n589, n588, \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q , 
        \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25_q , n600, n599, \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24_q , 
        \u_lcd_driver/r_lcd_rgb[5]~FF_frt_23_q , \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22_q , 
        \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21_q , \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q , 
        n613, n612, n611, n610, \u_lcd_driver/r_lcd_rgb[0]~FF_frt_19_q , 
        \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18_q , \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_q , 
        \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_q , \u_lcd_driver/r_lcd_dv~FF_frt_7_q , 
        \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q , \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2_q , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1_q , 
        \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_q , 
        n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, 
        n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, 
        n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, 
        n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, 
        n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, 
        n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, 
        n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, 
        n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, 
        n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, 
        n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, 
        n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, 
        n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, 
        n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, 
        n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, 
        n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, 
        n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, 
        n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, 
        n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, 
        n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, 
        n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, 
        n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, 
        n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, 
        n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, 
        n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, 
        n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, 
        n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, 
        n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, 
        n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, 
        n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, 
        n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, 
        n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, 
        n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, 
        n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, 
        n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, 
        n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, 
        n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, 
        n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, 
        n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, 
        n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, 
        n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, 
        n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, 
        n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, 
        n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, 
        n7381, n7383, n7399, n7400, n7401, n7402, n7403, n7404, 
        n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, 
        n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, 
        n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, 
        n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, 
        n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, 
        n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, 
        n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, 
        n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, 
        n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, 
        n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, 
        n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, 
        n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, 
        n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, 
        n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, 
        n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, 
        n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, 
        n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, 
        n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, 
        n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, 
        n7559, n7560, n7561;
    
    assign DdrCtrl_AID_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[31] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[30] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[29] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[28] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[27] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[26] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[9] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[8] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[5] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[4] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[3] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[2] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[1] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[2] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ABURST_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ABURST_0[0] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALOCK_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALOCK_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[15] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[14] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[13] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[12] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[11] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[10] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[9] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[8] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[7] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[6] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[5] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[4] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[3] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[2] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[1] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[0] = DdrCtrl_ALEN_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign cmos_ctl0 = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign cmos_ctl2 = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign cmos_ctl3 = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[4] = hdmi_txc_o[2] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[3] = hdmi_txc_o[2] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[1] = hdmi_txc_o[2] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign hdmi_txc_o[0] = hdmi_txc_o[2] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lcd_pwm = 1'b1 /* verific EFX_ATTRIBUTE_CELL_NAME=VCC */ ;
    assign lvds_tx0_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_LUT4 LUT__10591 (.I0(\u_axi4_ctrl/state[1] ), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(\u_axi4_ctrl/state[2] ), .O(DdrCtrl_AVALID_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__10591.LUTMASK = 16'h1414;
    EFX_FF \ResetShiftReg[0]~FF  (.D(\reduce_nand_9/n7 ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\ResetShiftReg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(128)
    defparam \ResetShiftReg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .CE_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .D_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_SYNC = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_VALUE = 1'b0;
    defparam \ResetShiftReg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[0]~FF  (.D(DdrInitDone), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(161)
    defparam \Axi0ResetReg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_rst_n~FF  (.D(\Axi0ResetReg[2] ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(r_hdmi_rst_n)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(456)
    defparam \r_hdmi_rst_n~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .SR_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_rst_n~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_rst_n~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_rst_n~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \rc_hdmi_tx~FF  (.D(rc_hdmi_tx), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(rc_hdmi_tx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \rc_hdmi_tx~FF .CLK_POLARITY = 1'b1;
    defparam \rc_hdmi_tx~FF .CE_POLARITY = 1'b1;
    defparam \rc_hdmi_tx~FF .SR_POLARITY = 1'b1;
    defparam \rc_hdmi_tx~FF .D_POLARITY = 1'b0;
    defparam \rc_hdmi_tx~FF .SR_SYNC = 1'b1;
    defparam \rc_hdmi_tx~FF .SR_VALUE = 1'b0;
    defparam \rc_hdmi_tx~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[0]~FF  (.D(n592_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx0_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[0]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[0]~FF  (.D(n603_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx1_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[0]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[0]~FF  (.D(n614_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx2_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[0]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[0]~FF  (.D(n3473), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ResetShiftReg[1]~FF  (.D(\ResetShiftReg[0] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\ResetShiftReg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(128)
    defparam \ResetShiftReg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .CE_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .D_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_SYNC = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_VALUE = 1'b0;
    defparam \ResetShiftReg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_CFG_RST_N~FF  (.D(\ResetShiftReg[1] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(DdrCtrl_CFG_RST_N)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(128)
    defparam \DdrCtrl_CFG_RST_N~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[1]~FF  (.D(\Axi0ResetReg[0] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(161)
    defparam \Axi0ResetReg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[2]~FF  (.D(\Axi0ResetReg[1] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(161)
    defparam \Axi0ResetReg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrInitDone~FF  (.D(1'b1), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(DdrInitDone)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \DdrInitDone~FF .CLK_POLARITY = 1'b1;
    defparam \DdrInitDone~FF .CE_POLARITY = 1'b0;
    defparam \DdrInitDone~FF .SR_POLARITY = 1'b0;
    defparam \DdrInitDone~FF .D_POLARITY = 1'b1;
    defparam \DdrInitDone~FF .SR_SYNC = 1'b0;
    defparam \DdrInitDone~FF .SR_VALUE = 1'b0;
    defparam \DdrInitDone~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_CFG_SEQ_START~FF  (.D(1'b1), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/equal_21/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(DdrCtrl_CFG_SEQ_START)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(186)
    defparam \DdrCtrl_CFG_SEQ_START~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_SEQ_START~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n92 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(186)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(150)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(150)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF  (.D(n176), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n91 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(186)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF  (.D(n3423), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF  (.D(n3421), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF  (.D(n3419), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF  (.D(n3417), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF  (.D(n3415), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF  (.D(n3413), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF  (.D(n3411), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF  (.D(n3409), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF  (.D(n3407), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF  (.D(n3405), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF  (.D(n3403), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF  (.D(n3401), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF  (.D(n3399), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF  (.D(n3397), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF  (.D(n3395), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF  (.D(n3393), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF  (.D(n3391), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF  (.D(n3389), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF  (.D(n3388), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n137 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(167)
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(167)
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n138 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n139 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n140 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n205 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[0]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[0]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[0]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[0]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n122 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n123 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n124 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n125 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n126 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n127 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n128 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n129 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n130 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n131 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n132 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n133 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n134 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n135 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n136 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(121)
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n500 ), 
           .CE(ceg_net552), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n509 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n567 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n570 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n573 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n576 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n579 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n581 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_capture_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(548)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .SR_VALUE = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_ack~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF  (.D(n197), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \cmos_sdat_OUT~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n495 ), .CE(ceg_net632), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(cmos_sdat_OUT)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \cmos_sdat_OUT~FF .CLK_POLARITY = 1'b1;
    defparam \cmos_sdat_OUT~FF .CE_POLARITY = 1'b1;
    defparam \cmos_sdat_OUT~FF .SR_POLARITY = 1'b0;
    defparam \cmos_sdat_OUT~FF .D_POLARITY = 1'b1;
    defparam \cmos_sdat_OUT~FF .SR_SYNC = 1'b0;
    defparam \cmos_sdat_OUT~FF .SR_VALUE = 1'b1;
    defparam \cmos_sdat_OUT~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(167)
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(167)
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(167)
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/current_state[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[1]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n204 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[1]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[1]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[1]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[1]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[2]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n203 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[2]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[2]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[2]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[2]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[2]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[3]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n202 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[3]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[3]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[3]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[3]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[3]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[4]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n201 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[4]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[4]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[4]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[4]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[4]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[5]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n200 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[5]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[5]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[5]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[5]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[5]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[6]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n199 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[6]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[6]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[6]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[6]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[6]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[6]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i2c_config_index[7]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n198 ), 
           .CE(\u_i2c_timing_ctrl_16reg_16bit/n846 ), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(\i2c_config_index[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(197)
    defparam \i2c_config_index[7]~FF .CLK_POLARITY = 1'b1;
    defparam \i2c_config_index[7]~FF .CE_POLARITY = 1'b1;
    defparam \i2c_config_index[7]~FF .SR_POLARITY = 1'b0;
    defparam \i2c_config_index[7]~FF .D_POLARITY = 1'b1;
    defparam \i2c_config_index[7]~FF .SR_SYNC = 1'b0;
    defparam \i2c_config_index[7]~FF .SR_VALUE = 1'b0;
    defparam \i2c_config_index[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n499 ), 
           .CE(ceg_net552), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n498 ), 
           .CE(ceg_net552), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n497 ), 
           .CE(ceg_net552), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n508 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n507 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n506 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n505 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n504 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n503 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF  (.D(\u_i2c_timing_ctrl_16reg_16bit/n502 ), 
           .CE(ceg_net664), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(497)
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF  (.D(n3382), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF  (.D(n3380), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF  (.D(n3378), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF  (.D(n3376), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF  (.D(n3374), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF  (.D(n3372), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF  (.D(n3370), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF  (.D(n3360), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF  (.D(n3358), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF  (.D(n3356), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF  (.D(n3354), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF  (.D(n3352), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF  (.D(n3350), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF  (.D(n3348), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF  (.D(n3346), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF  (.D(n3344), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF  (.D(n3342), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF  (.D(n3341), .CE(\u_i2c_timing_ctrl_16reg_16bit/n7 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(71)
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .SR_POLARITY = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .D_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .SR_SYNC = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .SR_VALUE = 1'b0;
    defparam \u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF  (.D(cmos_href), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_href_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF  (.D(cmos_data[0]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF  (.D(cmos_data[5]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n127 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF  (.D(cmos_data[4]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n160 ), 
           .CE(ceg_net158), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(128)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF  (.D(cmos_data[3]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF  (.D(1'b1), .CE(\u_CMOS_Capture_RAW_Gray/n171 ), 
           .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/frame_sync_flag )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(141)
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/frame_sync_flag~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF  (.D(cmos_data[2]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF  (.D(cmos_data[1]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF  (.D(cmos_data[7]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF  (.D(cmos_data[6]), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_data_r0[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_data_r0[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_href_r[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_href_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_href_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF  (.D(cmos_vsync), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n126 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n125 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n124 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n123 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n122 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n121 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n120 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n119 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n118 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n117 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n116 ), 
           .CE(ceg_net152), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/line_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(111)
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/line_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF  (.D(\u_CMOS_Capture_RAW_Gray/n159 ), 
           .CE(ceg_net158), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(128)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF  (.D(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(80)
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[9]~FF  (.D(\u_sensor_frame_count/n66 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[8]~FF  (.D(\u_sensor_frame_count/n67 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[7]~FF  (.D(\u_sensor_frame_count/n68 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[6]~FF  (.D(\u_sensor_frame_count/n69 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[5]~FF  (.D(\u_sensor_frame_count/n70 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[4]~FF  (.D(\u_sensor_frame_count/n71 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[1]~FF  (.D(\u_sensor_frame_count/n74 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[0]~FF  (.D(\u_sensor_frame_count/n141 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[3]~FF  (.D(\u_sensor_frame_count/n72 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[2]~FF  (.D(\u_sensor_frame_count/n73 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[0]~FF  (.D(\u_sensor_frame_count/n75 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[0]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[1] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[0]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[0]~FF .CE_POLARITY = 1'b0;
    defparam \LED[0]~FF .SR_POLARITY = 1'b0;
    defparam \LED[0]~FF .D_POLARITY = 1'b1;
    defparam \LED[0]~FF .SR_SYNC = 1'b0;
    defparam \LED[0]~FF .SR_VALUE = 1'b0;
    defparam \LED[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_vsync_r[0]~FF  (.D(cmos_vsync), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/cmos_vsync_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(53)
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[10]~FF  (.D(\u_sensor_frame_count/n65 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[11]~FF  (.D(\u_sensor_frame_count/n64 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[12]~FF  (.D(\u_sensor_frame_count/n63 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[13]~FF  (.D(\u_sensor_frame_count/n62 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[14]~FF  (.D(\u_sensor_frame_count/n61 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[15]~FF  (.D(\u_sensor_frame_count/n60 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[16]~FF  (.D(\u_sensor_frame_count/n59 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[17]~FF  (.D(\u_sensor_frame_count/n58 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[18]~FF  (.D(\u_sensor_frame_count/n57 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[19]~FF  (.D(\u_sensor_frame_count/n56 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[20]~FF  (.D(\u_sensor_frame_count/n55 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[21]~FF  (.D(\u_sensor_frame_count/n54 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[22]~FF  (.D(\u_sensor_frame_count/n53 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[23]~FF  (.D(\u_sensor_frame_count/n52 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[24]~FF  (.D(\u_sensor_frame_count/n51 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[25]~FF  (.D(\u_sensor_frame_count/n50 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[26]~FF  (.D(\u_sensor_frame_count/n49 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/delay_cnt[27]~FF  (.D(\u_sensor_frame_count/n48 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/delay_cnt[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(71)
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/delay_cnt[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[1]~FF  (.D(\u_sensor_frame_count/n140 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[2]~FF  (.D(\u_sensor_frame_count/n139 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[3]~FF  (.D(\u_sensor_frame_count/n138 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[4]~FF  (.D(\u_sensor_frame_count/n137 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[5]~FF  (.D(\u_sensor_frame_count/n136 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[6]~FF  (.D(\u_sensor_frame_count/n135 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[7]~FF  (.D(\u_sensor_frame_count/n134 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_fps_cnt[8]~FF  (.D(\u_sensor_frame_count/n133 ), 
           .CE(ceg_net200), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_sensor_frame_count/cmos_fps_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_fps_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[1]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[2] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[1]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[1]~FF .CE_POLARITY = 1'b0;
    defparam \LED[1]~FF .SR_POLARITY = 1'b0;
    defparam \LED[1]~FF .D_POLARITY = 1'b1;
    defparam \LED[1]~FF .SR_SYNC = 1'b0;
    defparam \LED[1]~FF .SR_VALUE = 1'b0;
    defparam \LED[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[2]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[3] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[2]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[2]~FF .CE_POLARITY = 1'b0;
    defparam \LED[2]~FF .SR_POLARITY = 1'b0;
    defparam \LED[2]~FF .D_POLARITY = 1'b1;
    defparam \LED[2]~FF .SR_SYNC = 1'b0;
    defparam \LED[2]~FF .SR_VALUE = 1'b0;
    defparam \LED[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[3]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[4] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[3]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[3]~FF .CE_POLARITY = 1'b0;
    defparam \LED[3]~FF .SR_POLARITY = 1'b0;
    defparam \LED[3]~FF .D_POLARITY = 1'b1;
    defparam \LED[3]~FF .SR_SYNC = 1'b0;
    defparam \LED[3]~FF .SR_VALUE = 1'b0;
    defparam \LED[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[4]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[5] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[4]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[4]~FF .CE_POLARITY = 1'b0;
    defparam \LED[4]~FF .SR_POLARITY = 1'b0;
    defparam \LED[4]~FF .D_POLARITY = 1'b1;
    defparam \LED[4]~FF .SR_SYNC = 1'b0;
    defparam \LED[4]~FF .SR_VALUE = 1'b0;
    defparam \LED[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[5]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[6] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[5]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[5]~FF .CE_POLARITY = 1'b0;
    defparam \LED[5]~FF .SR_POLARITY = 1'b0;
    defparam \LED[5]~FF .D_POLARITY = 1'b1;
    defparam \LED[5]~FF .SR_SYNC = 1'b0;
    defparam \LED[5]~FF .SR_VALUE = 1'b0;
    defparam \LED[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[6]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[7] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[6]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[6]~FF .CE_POLARITY = 1'b0;
    defparam \LED[6]~FF .SR_POLARITY = 1'b0;
    defparam \LED[6]~FF .D_POLARITY = 1'b1;
    defparam \LED[6]~FF .SR_SYNC = 1'b0;
    defparam \LED[6]~FF .SR_VALUE = 1'b0;
    defparam \LED[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \LED[7]~FF  (.D(\u_sensor_frame_count/cmos_fps_cnt[8] ), .CE(\u_sensor_frame_count/n110 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(LED[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(94)
    defparam \LED[7]~FF .CLK_POLARITY = 1'b1;
    defparam \LED[7]~FF .CE_POLARITY = 1'b0;
    defparam \LED[7]~FF .SR_POLARITY = 1'b0;
    defparam \LED[7]~FF .D_POLARITY = 1'b1;
    defparam \LED[7]~FF .SR_SYNC = 1'b0;
    defparam \LED[7]~FF .SR_VALUE = 1'b0;
    defparam \LED[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_sensor_frame_count/cmos_vsync_r[1]~FF  (.D(\u_sensor_frame_count/cmos_vsync_r[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_sensor_frame_count/cmos_vsync_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(53)
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_sensor_frame_count/cmos_vsync_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(499)
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF  (.D(1'b0), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(499)
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF  (.D(1'b0), .CE(1'b1), 
           .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(492)
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(721)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF  (.D(n2799), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF  (.D(n2801), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/waddr[0] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), .CLK(\cmos_pclk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/waddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF  (.D(n2803), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF  (.D(n681), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \empty~FF  (.D(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CE(ceg_net219), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(empty)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1090)
    defparam \empty~FF .CLK_POLARITY = 1'b1;
    defparam \empty~FF .CE_POLARITY = 1'b0;
    defparam \empty~FF .SR_POLARITY = 1'b1;
    defparam \empty~FF .D_POLARITY = 1'b0;
    defparam \empty~FF .SR_SYNC = 1'b0;
    defparam \empty~FF .SR_VALUE = 1'b1;
    defparam \empty~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF  (.D(n2805), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF  (.D(n2807), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/raddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF  (.D(n2809), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF  (.D(n2811), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF  (.D(n703), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF  (.D(n2797), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF  (.D(n2795), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF  (.D(n2793), .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
           .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/waddr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/waddr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF  (.D(n2792), 
           .CE(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), .CLK(\cmos_pclk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1273)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF  (.D(n715), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF  (.D(n2776), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF  (.D(n2774), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF  (.D(n2772), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF  (.D(n2770), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF  (.D(n2768), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF  (.D(n2766), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF  (.D(n2764), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF  (.D(n2762), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF  (.D(n2760), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF  (.D(n2758), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF  (.D(n2756), .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/raddr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/raddr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF  (.D(n2755), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[1] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[2] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[3] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[4] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[5] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[6] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[7] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[8] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[9] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[10] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[11] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] ), 
           .CE(\u_afifo_buf/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1284)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[13] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1339)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[12] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1351)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[13] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[13] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2  (.D(n7112), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true", INIT_VALUE=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1  (.D(n6311), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true", INIT_VALUE=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1 .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1 .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1 .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1 .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1 .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1 .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF  (.D(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[0] ), 
           .CE(1'b1), .CLK(\cmos_pclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(492)
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[0]~FF  (.D(\u_scaler_gray/vs_cnt[0] ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tvsync_o~FF  (.D(\u_scaler_gray/n150 ), .CE(ceg_net229), .CLK(\Axi_Clk~O ), 
           .SR(\Axi0ResetReg[2] ), .Q(tvsync_o)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(123)
    defparam \tvsync_o~FF .CLK_POLARITY = 1'b1;
    defparam \tvsync_o~FF .CE_POLARITY = 1'b0;
    defparam \tvsync_o~FF .SR_POLARITY = 1'b0;
    defparam \tvsync_o~FF .D_POLARITY = 1'b0;
    defparam \tvsync_o~FF .SR_SYNC = 1'b0;
    defparam \tvsync_o~FF .SR_VALUE = 1'b0;
    defparam \tvsync_o~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] ), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/tvalid_o_r~FF  (.D(tvalid_o), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\u_scaler_gray/tvalid_o_r )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(97)
    defparam \u_scaler_gray/tvalid_o_r~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid_o_r~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid_o_r~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid_o_r~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid_o_r~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/tvalid_o_r~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/tvalid_o_r~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/w_addra[0] ), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n432 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(176)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n2156 ), 
           .CE(ceg_net526), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(176)
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[0]~FF  (.D(\u_scaler_gray/destx[0] ), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[0]~FF  (.D(\u_scaler_gray/desty[0] ), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/desty[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n903 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n903 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0] ), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF  (.D(n904), .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF  (.D(n2543), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF  (.D(n2541), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF  (.D(n2539), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF  (.D(n2527), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF  (.D(n2522), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF  (.D(n2498), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF  (.D(n2496), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF  (.D(n2494), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF  (.D(n2492), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF  (.D(n2490), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF  (.D(n2488), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF  (.D(n2486), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF  (.D(n2484), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF  (.D(n2483), 
           .CE(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast ), .CLK(\Axi_Clk~O ), 
           .SR(\u_scaler_gray/u0_data_stream_ctr/n1703 ), .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(81)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF  (.D(n911), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF  (.D(n2402), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF  (.D(n2400), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF  (.D(n2398), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF  (.D(n2396), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF  (.D(n2394), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF  (.D(n2392), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF  (.D(n2382), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF  (.D(n2380), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF  (.D(n2378), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF  (.D(n2376), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF  (.D(n2374), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF  (.D(n2372), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF  (.D(n2370), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF  (.D(n2369), .CE(n197_2), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1704 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_addra[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(94)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_addra[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n431 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(176)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n430 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(176)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_st[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n2073 ), 
           .CE(ceg_net526), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(176)
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/delay_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[1]~FF  (.D(n916), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[2]~FF  (.D(n2352), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[3]~FF  (.D(n2346), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[4]~FF  (.D(n2343), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[5]~FF  (.D(n2338), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[6]~FF  (.D(n2336), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[7]~FF  (.D(n2334), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[8]~FF  (.D(n2330), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[9]~FF  (.D(n2328), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[9]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[10]~FF  (.D(n2326), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[10]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[11]~FF  (.D(n2324), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[11]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[12]~FF  (.D(n2322), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[12]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[13]~FF  (.D(n2320), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[13]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[14]~FF  (.D(n2315), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[14]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/destx[15]~FF  (.D(n2314), .CE(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1712 ), 
           .Q(\u_scaler_gray/destx[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(195)
    defparam \u_scaler_gray/destx[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[15]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/destx[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/destx[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/destx[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/destx[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[1]~FF  (.D(n934), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[2]~FF  (.D(n2312), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[3]~FF  (.D(n2304), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[4]~FF  (.D(n2302), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[5]~FF  (.D(n2300), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[6]~FF  (.D(n2298), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[7]~FF  (.D(n2296), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[8]~FF  (.D(n2291), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[9]~FF  (.D(n2234), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[10]~FF  (.D(n2232), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[11]~FF  (.D(n2230), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[12]~FF  (.D(n2228), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[13]~FF  (.D(n2226), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[14]~FF  (.D(n2224), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/desty[15]~FF  (.D(n2187), .CE(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
           .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1713 ), 
           .Q(\u_scaler_gray/desty[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(214)
    defparam \u_scaler_gray/desty[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/desty[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/desty[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/desty[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1196 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1161 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1160 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1159 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n885 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n884 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n883 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n882 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n881 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n880 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n879 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1179 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1178 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1177 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1176 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF  (.D(\u_scaler_gray/srcx_int[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF  (.D(\u_scaler_gray/srcx_int[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF  (.D(\u_scaler_gray/srcx_int[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF  (.D(\u_scaler_gray/srcx_int[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF  (.D(\u_scaler_gray/srcx_int[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF  (.D(\u_scaler_gray/srcx_int[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF  (.D(\u_scaler_gray/srcx_int[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1196 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1195 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1194 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1193 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1179 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1212 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1211 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/n1210 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(247)
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/tvalid~FF  (.D(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/tvalid )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(265)
    defparam \u_scaler_gray/tvalid~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/tvalid~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/tvalid~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/tvalid~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF  (.D(n735), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF  (.D(n2692), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF  (.D(n2690), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF  (.D(n2686), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF  (.D(n2683), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF  (.D(n2681), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF  (.D(n2679), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF  (.D(n2597), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF  (.D(n2595), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF  (.D(n2593), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF  (.D(n2591), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF  (.D(n2589), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF  (.D(n2587), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF  (.D(n2585), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF  (.D(n2584), 
           .CE(n197_2), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u0_data_stream_ctr/n1702 ), 
           .Q(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(63)
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[1]~FF  (.D(\u_scaler_gray/n129 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[2]~FF  (.D(\u_scaler_gray/n128 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[3]~FF  (.D(\u_scaler_gray/n127 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[4]~FF  (.D(\u_scaler_gray/n126 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[5]~FF  (.D(\u_scaler_gray/n125 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[6]~FF  (.D(\u_scaler_gray/n124 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[7]~FF  (.D(\u_scaler_gray/n123 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[8]~FF  (.D(\u_scaler_gray/n122 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[9]~FF  (.D(\u_scaler_gray/n121 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[10]~FF  (.D(\u_scaler_gray/n120 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[11]~FF  (.D(\u_scaler_gray/n119 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[12]~FF  (.D(\u_scaler_gray/n118 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[12]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[13]~FF  (.D(\u_scaler_gray/n117 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[13]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[14]~FF  (.D(\u_scaler_gray/n116 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[14]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/vs_cnt[15]~FF  (.D(\u_scaler_gray/n115 ), .CE(ceg_net226), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/vs_cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(111)
    defparam \u_scaler_gray/vs_cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[15]~FF .CE_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/vs_cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/vs_cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \u_scaler_gray/vs_cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/vs_cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n462 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ASIZE_0[2]~FF  (.D(1'b1), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(DdrCtrl_ALEN_0[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \DdrCtrl_ASIZE_0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ASIZE_0[2]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ASIZE_0[2]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ASIZE_0[2]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ASIZE_0[2]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_ASIZE_0[2]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ASIZE_0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF  (.D(n2169), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF  (.D(n2166), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF  (.D(n2164), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF  (.D(n2162), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF  (.D(n2160), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF  (.D(n2158), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF  (.D(n2155), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF  (.D(n2153), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF  (.D(n2151), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF  (.D(n2147), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF  (.D(n2144), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF  (.D(n2142), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF  (.D(n2140), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF  (.D(n2138), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF  (.D(n2136), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF  (.D(n2133), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF  (.D(n2132), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF  (.D(n1534), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF  (.D(n2126), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF  (.D(n2122), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF  (.D(n2119), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF  (.D(n2115), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF  (.D(n2112), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF  (.D(n2109), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF  (.D(n2107), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF  (.D(n2066), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF  (.D(n2064), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF  (.D(n2062), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF  (.D(n2060), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF  (.D(n2058), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF  (.D(n2056), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF  (.D(n2054), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF  (.D(n1769), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF  (.D(n1713), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF  (.D(n1692), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF  (.D(n1690), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF  (.D(n1688), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF  (.D(n1686), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF  (.D(n1684), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF  (.D(n1682), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF  (.D(n1680), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF  (.D(n1678), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF  (.D(n1676), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF  (.D(n1671), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(63)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__10592 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/wdata_cnt_dly[4] ), 
            .O(n7037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10592.LUTMASK = 16'h0001;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n335 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcx_fix[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n334 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcx_fix[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n333 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcx_fix[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcx_fix[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n332 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n331 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n330 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n329 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n328 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n327 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n326 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n325 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[8]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n324 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n323 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n322 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n321 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[12]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n320 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[13]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n319 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[14]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n318 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcx_int[15]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n317 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcx_int[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(72)
    defparam \u_scaler_gray/srcx_int[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcx_int[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcx_int[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcx_int[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n461 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n460 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n459 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n458 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n457 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n456 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n455 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n454 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n453 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n452 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n451 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/srcy_fix[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/srcy_fix[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n450 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n449 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n448 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n447 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n446 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n445 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n444 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n443 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[8]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n442 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n441 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n440 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n439 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[12]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n438 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[13]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n437 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[14]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n436 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/srcy_int[15]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n435 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/srcy_int[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(81)
    defparam \u_scaler_gray/srcy_int[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/srcy_int[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/srcy_int[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/srcy_int[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF  (.D(\u_scaler_gray/destx[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF  (.D(\u_scaler_gray/destx[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF  (.D(n1536), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF  (.D(n1515), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF  (.D(n1513), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF  (.D(n1511), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF  (.D(n1509), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF  (.D(n1507), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF  (.D(n1505), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF  (.D(n1503), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF  (.D(n1501), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF  (.D(n1499), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF  (.D(n1497), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF  (.D(n1495), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF  (.D(n1480), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF  (.D(n1478), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF  (.D(n1476), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF  (.D(n1475), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(26)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcy_fix[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcx_fix[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(26)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcx_fix[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(26)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/srcx_fix[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(26)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .D_POLARITY = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF  (.D(n1739), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF  (.D(n1908), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n344 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[0]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[0]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[0]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[0]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[0]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[0]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[0]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF  (.D(\u_scaler_gray/tvalid ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_GBUFCE CLKBUF__3 (.CE(1'b1), .I(cmos_pclk), .O(\cmos_pclk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__3.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__2 (.CE(1'b1), .I(hdmi_clk2x_i), .O(\hdmi_clk2x_i~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__2.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(hdmi_clk1x_i), .O(\hdmi_clk1x_i~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF  (.D(n1101), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF  (.D(n1099), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF  (.D(n1097), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF  (.D(n1095), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF  (.D(n1093), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF  (.D(n1091), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF  (.D(n1089), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF  (.D(n1087), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF  (.D(n1085), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF  (.D(n1083), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF  (.D(n1081), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF  (.D(n1079), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF  (.D(n1077), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF  (.D(n1075), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF  (.D(n1073), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF  (.D(n1071), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF  (.D(n1069), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF  (.D(n1067), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF  (.D(n1065), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF  (.D(n1066), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF  (.D(n1048), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF  (.D(n1046), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF  (.D(n1044), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF  (.D(n1042), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF  (.D(n1040), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF  (.D(n1038), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF  (.D(n1036), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF  (.D(n1034), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF  (.D(n1032), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF  (.D(n1030), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF  (.D(n1028), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF  (.D(n1026), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF  (.D(n1024), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF  (.D(n1022), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF  (.D(n1020), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF  (.D(n1018), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF  (.D(n1016), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF  (.D(n1014), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF  (.D(n1012), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF  (.D(n1013), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(43)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF  (.D(n958), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF  (.D(n956), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF  (.D(n954), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF  (.D(n952), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF  (.D(n950), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF  (.D(n948), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF  (.D(n946), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF  (.D(n944), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF  (.D(n942), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF  (.D(n940), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF  (.D(n941), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(48)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n343 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n342 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n341 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n340 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n339 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n338 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n337 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n336 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n335 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(60)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[1]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[1]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[1]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[2]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[2]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[2]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[3]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[3]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[3]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[4]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[4]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[4]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[4]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[5]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[5]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[5]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[5]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[5]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[5]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[5]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[6]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[6]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[6]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[6]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[6]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tdata_o[7]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 ), 
           .Q(\tdata_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(65)
    defparam \tdata_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \tdata_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \tdata_o[7]~FF .SR_POLARITY = 1'b1;
    defparam \tdata_o[7]~FF .D_POLARITY = 1'b1;
    defparam \tdata_o[7]~FF .SR_SYNC = 1'b1;
    defparam \tdata_o[7]~FF .SR_VALUE = 1'b1;
    defparam \tdata_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .D_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .SR_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .SR_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tvalid_o~FF  (.D(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/tvalid_d[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(tvalid_o)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(70)
    defparam \tvalid_o~FF .CLK_POLARITY = 1'b1;
    defparam \tvalid_o~FF .CE_POLARITY = 1'b1;
    defparam \tvalid_o~FF .SR_POLARITY = 1'b1;
    defparam \tvalid_o~FF .D_POLARITY = 1'b1;
    defparam \tvalid_o~FF .SR_SYNC = 1'b1;
    defparam \tvalid_o~FF .SR_VALUE = 1'b0;
    defparam \tvalid_o~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(Axi_Clk), .O(\Axi_Clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_52/add_2/i2  (.I0(n3336), .I1(1'b1), 
            .CI(1'b0), .CO(n7579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(79)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_52/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_52/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_50/add_2/i2  (.I0(n3336), .I1(1'b1), 
            .CI(1'b0), .CO(n7578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_50/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_50/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__u_rgb2dvi/enc_2/sub_50/add_2/i1  (.I0(1'b0), .I1(1'b0), 
            .CI(n7577), .O(n3336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \AUX_ADD_CO__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_2/sub_50/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n7576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_2/sub_50/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_79/add_2/i2  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n7575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(93)
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_79/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_rgb2dvi/enc_0/sub_79/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n7574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n7572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n7571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n7570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n7569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n7568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n7567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20  (.I0(1'b0), 
            .I1(1'b0), .CI(n7566), .O(n1066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20  (.I0(1'b0), 
            .I1(1'b0), .CI(n7565), .O(n1013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21  (.I0(1'b0), 
            .I1(1'b0), .CI(n7564), .O(n941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n7563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \AUX_ADD_CI__u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n7562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[0]~FF  (.D(tvsync_o), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_index[1]~FF  (.D(\u_axi4_ctrl/n316 ), .CE(\u_axi4_ctrl/equal_38/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(177)
    defparam \u_axi4_ctrl/wframe_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[0]~FF  (.D(lcd_vs), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_index[0]~FF  (.D(\u_axi4_ctrl/n317 ), .CE(\u_axi4_ctrl/equal_38/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(177)
    defparam \u_axi4_ctrl/wframe_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF  (.D(n741), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_index[0]~FF  (.D(\u_axi4_ctrl/n336 ), .CE(\u_axi4_ctrl/equal_47/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(197)
    defparam \u_axi4_ctrl/rframe_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/state[0]~FF  (.D(\u_axi4_ctrl/n389 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(268)
    defparam \u_axi4_ctrl/state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/state[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[1]~FF  (.D(\u_axi4_ctrl/wframe_vsync_dly[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ATYPE_0~FF  (.D(1'b1), .CE(\u_axi4_ctrl/n405 ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/n1476 ), .Q(DdrCtrl_ATYPE_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(283)
    defparam \DdrCtrl_ATYPE_0~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ATYPE_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[3]~FF  (.D(\u_axi4_ctrl/wframe_vsync_dly[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF  (.D(n2269), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF  (.D(n2271), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[0]~FF  (.D(\u_axi4_ctrl/wdata_cnt_dly[0] ), 
           .CE(\u_axi4_ctrl/n363 ), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), 
           .Q(\u_axi4_ctrl/wdata_cnt_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[1]~FF  (.D(\u_axi4_ctrl/n1544 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[0]~FF  (.D(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
           .CE(\u_axi4_ctrl/n379 ), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), 
           .Q(\u_axi4_ctrl/rdata_cnt_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[3]~FF  (.D(\u_axi4_ctrl/rframe_vsync_dly[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[2]~FF  (.D(\u_axi4_ctrl/rframe_vsync_dly[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wenb~FF  (.D(\u_axi4_ctrl/n379 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rfifo_wenb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(434)
    defparam \u_axi4_ctrl/rfifo_wenb~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[1]~FF  (.D(\u_axi4_ctrl/rframe_vsync_dly[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[0]~FF  (.D(DdrCtrl_RDATA_0[0]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[2]~FF  (.D(\u_axi4_ctrl/wframe_vsync_dly[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(79)
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF  (.D(n739), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wfifo_empty~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CE(ceg_net289), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/wfifo_empty )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1090)
    defparam \u_axi4_ctrl/wfifo_empty~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_empty~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_empty~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF  (.D(n743), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF  (.D(n672), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF  (.D(n683), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF  (.D(n712), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF  (.D(n718), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF  (.D(n723), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF  (.D(n737), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF  (.D(n745), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF  (.D(n2349), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF  (.D(n670), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF  (.D(n668), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF  (.D(n666), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF  (.D(n664), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF  (.D(n662), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF  (.D(n660), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF  (.D(n659), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_empty~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CE(ceg_net296), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/rfifo_empty )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1090)
    defparam \u_axi4_ctrl/rfifo_empty~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_empty~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_empty~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF  (.D(n2512), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF  (.D(n2510), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF  (.D(n555), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF  (.D(n553), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF  (.D(n551), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF  (.D(n549), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF  (.D(n547), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF  (.D(n546), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF  (.D(n2517), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF  (.D(n544), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF  (.D(n542), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF  (.D(n540), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF  (.D(n538), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF  (.D(n536), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF  (.D(n534), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF  (.D(n524), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF  (.D(n479), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF  (.D(n466), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF  (.D(n464), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF  (.D(n457), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\hdmi_clk1x_i~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_index[1]~FF  (.D(\u_axi4_ctrl/n335 ), .CE(\u_axi4_ctrl/equal_47/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(197)
    defparam \u_axi4_ctrl/rframe_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/state[1]~FF  (.D(\u_axi4_ctrl/n1610 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1617 ), .Q(\u_axi4_ctrl/state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(268)
    defparam \u_axi4_ctrl/state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/state[2]~FF  (.D(\u_axi4_ctrl/n387 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(268)
    defparam \u_axi4_ctrl/state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/state[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[10]~FF  (.D(\u_axi4_ctrl/awaddr[10] ), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[11]~FF  (.D(n2149), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[12]~FF  (.D(n802), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[13]~FF  (.D(n800), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[14]~FF  (.D(n798), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[15]~FF  (.D(n796), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[16]~FF  (.D(n794), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[17]~FF  (.D(n792), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[18]~FF  (.D(n790), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[19]~FF  (.D(n788), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[20]~FF  (.D(n786), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[21]~FF  (.D(n784), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[22]~FF  (.D(n782), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[23]~FF  (.D(n781), .CE(\u_axi4_ctrl/n369 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1469 ), .Q(\u_axi4_ctrl/awaddr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(301)
    defparam \u_axi4_ctrl/awaddr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[10]~FF  (.D(\u_axi4_ctrl/araddr[10] ), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[11]~FF  (.D(n2124), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[12]~FF  (.D(n2188), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[13]~FF  (.D(n779), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[14]~FF  (.D(n777), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[15]~FF  (.D(n775), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[16]~FF  (.D(n773), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[17]~FF  (.D(n771), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[18]~FF  (.D(n769), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[19]~FF  (.D(n754), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[20]~FF  (.D(n752), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[21]~FF  (.D(n750), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[22]~FF  (.D(n748), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[23]~FF  (.D(n747), .CE(\u_axi4_ctrl/n381 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1478 ), .Q(\u_axi4_ctrl/araddr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(319)
    defparam \u_axi4_ctrl/araddr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[10]~FF  (.D(\u_axi4_ctrl/n697 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[10]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[10]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[10]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[11]~FF  (.D(\u_axi4_ctrl/n696 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[11]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[11]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[11]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[12]~FF  (.D(\u_axi4_ctrl/n695 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[12]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[12]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[12]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[13]~FF  (.D(\u_axi4_ctrl/n694 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[13]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[13]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[13]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[14]~FF  (.D(\u_axi4_ctrl/n693 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[14]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[14]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[14]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[15]~FF  (.D(\u_axi4_ctrl/n692 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[15]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[15]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[16]~FF  (.D(\u_axi4_ctrl/n691 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[16]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[16]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[16]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[17]~FF  (.D(\u_axi4_ctrl/n690 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[17]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[17]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[17]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[18]~FF  (.D(\u_axi4_ctrl/n689 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[18]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[18]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[18]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[19]~FF  (.D(\u_axi4_ctrl/n688 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[19]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[19]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[19]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[20]~FF  (.D(\u_axi4_ctrl/n687 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[20]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[20]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[20]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[21]~FF  (.D(\u_axi4_ctrl/n686 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[21]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[21]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[21]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[22]~FF  (.D(\u_axi4_ctrl/n685 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[22]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[22]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[22]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[23]~FF  (.D(\u_axi4_ctrl/n684 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[23]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[23]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[23]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[24]~FF  (.D(\u_axi4_ctrl/n683 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[24]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[24]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[24]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[25]~FF  (.D(\u_axi4_ctrl/n682 ), .CE(ceg_net401), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(334)
    defparam \DdrCtrl_AADDR_0[25]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[25]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[25]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[1]~FF  (.D(\u_axi4_ctrl/n1499 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[2]~FF  (.D(\u_axi4_ctrl/n1504 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[3]~FF  (.D(\u_axi4_ctrl/n1509 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[4]~FF  (.D(\u_axi4_ctrl/n1514 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[5]~FF  (.D(\u_axi4_ctrl/n1519 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[6]~FF  (.D(\u_axi4_ctrl/n1524 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[7]~FF  (.D(\u_axi4_ctrl/n1529 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[8]~FF  (.D(\u_axi4_ctrl/n1534 ), .CE(\u_axi4_ctrl/n363 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(349)
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[2]~FF  (.D(\u_axi4_ctrl/n1549 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[3]~FF  (.D(\u_axi4_ctrl/n1554 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[4]~FF  (.D(\u_axi4_ctrl/n1559 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[5]~FF  (.D(\u_axi4_ctrl/n1564 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[6]~FF  (.D(\u_axi4_ctrl/n1569 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[7]~FF  (.D(\u_axi4_ctrl/n1574 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[8]~FF  (.D(\u_axi4_ctrl/n1579 ), .CE(\u_axi4_ctrl/n379 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(400)
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[1]~FF  (.D(DdrCtrl_RDATA_0[1]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[2]~FF  (.D(DdrCtrl_RDATA_0[2]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[3]~FF  (.D(DdrCtrl_RDATA_0[3]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[4]~FF  (.D(DdrCtrl_RDATA_0[4]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[5]~FF  (.D(DdrCtrl_RDATA_0[5]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[6]~FF  (.D(DdrCtrl_RDATA_0[6]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[7]~FF  (.D(DdrCtrl_RDATA_0[7]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[8]~FF  (.D(DdrCtrl_RDATA_0[8]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[9]~FF  (.D(DdrCtrl_RDATA_0[9]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[10]~FF  (.D(DdrCtrl_RDATA_0[10]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[11]~FF  (.D(DdrCtrl_RDATA_0[11]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[12]~FF  (.D(DdrCtrl_RDATA_0[12]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[13]~FF  (.D(DdrCtrl_RDATA_0[13]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[14]~FF  (.D(DdrCtrl_RDATA_0[14]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[15]~FF  (.D(DdrCtrl_RDATA_0[15]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[16]~FF  (.D(DdrCtrl_RDATA_0[16]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[17]~FF  (.D(DdrCtrl_RDATA_0[17]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[18]~FF  (.D(DdrCtrl_RDATA_0[18]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[19]~FF  (.D(DdrCtrl_RDATA_0[19]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[20]~FF  (.D(DdrCtrl_RDATA_0[20]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[21]~FF  (.D(DdrCtrl_RDATA_0[21]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[22]~FF  (.D(DdrCtrl_RDATA_0[22]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[23]~FF  (.D(DdrCtrl_RDATA_0[23]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[24]~FF  (.D(DdrCtrl_RDATA_0[24]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[25]~FF  (.D(DdrCtrl_RDATA_0[25]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[26]~FF  (.D(DdrCtrl_RDATA_0[26]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[27]~FF  (.D(DdrCtrl_RDATA_0[27]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[28]~FF  (.D(DdrCtrl_RDATA_0[28]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[29]~FF  (.D(DdrCtrl_RDATA_0[29]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[30]~FF  (.D(DdrCtrl_RDATA_0[30]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[31]~FF  (.D(DdrCtrl_RDATA_0[31]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[32]~FF  (.D(DdrCtrl_RDATA_0[32]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[33]~FF  (.D(DdrCtrl_RDATA_0[33]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[34]~FF  (.D(DdrCtrl_RDATA_0[34]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[35]~FF  (.D(DdrCtrl_RDATA_0[35]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[36]~FF  (.D(DdrCtrl_RDATA_0[36]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[37]~FF  (.D(DdrCtrl_RDATA_0[37]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[38]~FF  (.D(DdrCtrl_RDATA_0[38]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[39]~FF  (.D(DdrCtrl_RDATA_0[39]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[40]~FF  (.D(DdrCtrl_RDATA_0[40]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[41]~FF  (.D(DdrCtrl_RDATA_0[41]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[42]~FF  (.D(DdrCtrl_RDATA_0[42]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[43]~FF  (.D(DdrCtrl_RDATA_0[43]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[44]~FF  (.D(DdrCtrl_RDATA_0[44]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[45]~FF  (.D(DdrCtrl_RDATA_0[45]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[46]~FF  (.D(DdrCtrl_RDATA_0[46]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[47]~FF  (.D(DdrCtrl_RDATA_0[47]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[48]~FF  (.D(DdrCtrl_RDATA_0[48]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[49]~FF  (.D(DdrCtrl_RDATA_0[49]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[50]~FF  (.D(DdrCtrl_RDATA_0[50]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[51]~FF  (.D(DdrCtrl_RDATA_0[51]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[52]~FF  (.D(DdrCtrl_RDATA_0[52]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[53]~FF  (.D(DdrCtrl_RDATA_0[53]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[54]~FF  (.D(DdrCtrl_RDATA_0[54]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[55]~FF  (.D(DdrCtrl_RDATA_0[55]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[56]~FF  (.D(DdrCtrl_RDATA_0[56]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[57]~FF  (.D(DdrCtrl_RDATA_0[57]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[58]~FF  (.D(DdrCtrl_RDATA_0[58]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[59]~FF  (.D(DdrCtrl_RDATA_0[59]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[60]~FF  (.D(DdrCtrl_RDATA_0[60]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[61]~FF  (.D(DdrCtrl_RDATA_0[61]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[62]~FF  (.D(DdrCtrl_RDATA_0[62]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[63]~FF  (.D(DdrCtrl_RDATA_0[63]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[64]~FF  (.D(DdrCtrl_RDATA_0[64]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[65]~FF  (.D(DdrCtrl_RDATA_0[65]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[66]~FF  (.D(DdrCtrl_RDATA_0[66]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[67]~FF  (.D(DdrCtrl_RDATA_0[67]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[68]~FF  (.D(DdrCtrl_RDATA_0[68]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[69]~FF  (.D(DdrCtrl_RDATA_0[69]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[70]~FF  (.D(DdrCtrl_RDATA_0[70]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[71]~FF  (.D(DdrCtrl_RDATA_0[71]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[72]~FF  (.D(DdrCtrl_RDATA_0[72]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[73]~FF  (.D(DdrCtrl_RDATA_0[73]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[74]~FF  (.D(DdrCtrl_RDATA_0[74]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[75]~FF  (.D(DdrCtrl_RDATA_0[75]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[76]~FF  (.D(DdrCtrl_RDATA_0[76]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[77]~FF  (.D(DdrCtrl_RDATA_0[77]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[78]~FF  (.D(DdrCtrl_RDATA_0[78]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[79]~FF  (.D(DdrCtrl_RDATA_0[79]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[80]~FF  (.D(DdrCtrl_RDATA_0[80]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[81]~FF  (.D(DdrCtrl_RDATA_0[81]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[82]~FF  (.D(DdrCtrl_RDATA_0[82]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[83]~FF  (.D(DdrCtrl_RDATA_0[83]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[84]~FF  (.D(DdrCtrl_RDATA_0[84]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[85]~FF  (.D(DdrCtrl_RDATA_0[85]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[86]~FF  (.D(DdrCtrl_RDATA_0[86]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[87]~FF  (.D(DdrCtrl_RDATA_0[87]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[88]~FF  (.D(DdrCtrl_RDATA_0[88]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[89]~FF  (.D(DdrCtrl_RDATA_0[89]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[90]~FF  (.D(DdrCtrl_RDATA_0[90]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[91]~FF  (.D(DdrCtrl_RDATA_0[91]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[92]~FF  (.D(DdrCtrl_RDATA_0[92]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[93]~FF  (.D(DdrCtrl_RDATA_0[93]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[94]~FF  (.D(DdrCtrl_RDATA_0[94]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[95]~FF  (.D(DdrCtrl_RDATA_0[95]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[96]~FF  (.D(DdrCtrl_RDATA_0[96]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[97]~FF  (.D(DdrCtrl_RDATA_0[97]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[98]~FF  (.D(DdrCtrl_RDATA_0[98]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[99]~FF  (.D(DdrCtrl_RDATA_0[99]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[100]~FF  (.D(DdrCtrl_RDATA_0[100]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[101]~FF  (.D(DdrCtrl_RDATA_0[101]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[102]~FF  (.D(DdrCtrl_RDATA_0[102]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[103]~FF  (.D(DdrCtrl_RDATA_0[103]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[104]~FF  (.D(DdrCtrl_RDATA_0[104]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[105]~FF  (.D(DdrCtrl_RDATA_0[105]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[106]~FF  (.D(DdrCtrl_RDATA_0[106]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[107]~FF  (.D(DdrCtrl_RDATA_0[107]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[108]~FF  (.D(DdrCtrl_RDATA_0[108]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[109]~FF  (.D(DdrCtrl_RDATA_0[109]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[110]~FF  (.D(DdrCtrl_RDATA_0[110]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[111]~FF  (.D(DdrCtrl_RDATA_0[111]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[112]~FF  (.D(DdrCtrl_RDATA_0[112]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[113]~FF  (.D(DdrCtrl_RDATA_0[113]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[114]~FF  (.D(DdrCtrl_RDATA_0[114]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[115]~FF  (.D(DdrCtrl_RDATA_0[115]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[116]~FF  (.D(DdrCtrl_RDATA_0[116]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[117]~FF  (.D(DdrCtrl_RDATA_0[117]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[118]~FF  (.D(DdrCtrl_RDATA_0[118]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[119]~FF  (.D(DdrCtrl_RDATA_0[119]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[120]~FF  (.D(DdrCtrl_RDATA_0[120]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[121]~FF  (.D(DdrCtrl_RDATA_0[121]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[122]~FF  (.D(DdrCtrl_RDATA_0[122]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[123]~FF  (.D(DdrCtrl_RDATA_0[123]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[124]~FF  (.D(DdrCtrl_RDATA_0[124]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[125]~FF  (.D(DdrCtrl_RDATA_0[125]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[126]~FF  (.D(DdrCtrl_RDATA_0[126]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[127]~FF  (.D(DdrCtrl_RDATA_0[127]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(439)
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[0]~FF  (.D(\u_lcd_driver/n83 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_hs~FF  (.D(\u_lcd_driver/n35 ), .CE(r_hdmi_rst_n), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(lcd_hs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \lcd_hs~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_hs~FF .CE_POLARITY = 1'b1;
    defparam \lcd_hs~FF .SR_POLARITY = 1'b1;
    defparam \lcd_hs~FF .D_POLARITY = 1'b0;
    defparam \lcd_hs~FF .SR_SYNC = 1'b1;
    defparam \lcd_hs~FF .SR_VALUE = 1'b0;
    defparam \lcd_hs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_vs~FF  (.D(\u_lcd_driver/n97 ), .CE(r_hdmi_rst_n), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(lcd_vs)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \lcd_vs~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_vs~FF .CE_POLARITY = 1'b1;
    defparam \lcd_vs~FF .SR_POLARITY = 1'b1;
    defparam \lcd_vs~FF .D_POLARITY = 1'b0;
    defparam \lcd_vs~FF .SR_SYNC = 1'b1;
    defparam \lcd_vs~FF .SR_VALUE = 1'b0;
    defparam \lcd_vs~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \lcd_de~FF  (.D(\u_lcd_driver/n125 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(lcd_de)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \lcd_de~FF .CLK_POLARITY = 1'b1;
    defparam \lcd_de~FF .CE_POLARITY = 1'b1;
    defparam \lcd_de~FF .SR_POLARITY = 1'b1;
    defparam \lcd_de~FF .D_POLARITY = 1'b1;
    defparam \lcd_de~FF .SR_SYNC = 1'b1;
    defparam \lcd_de~FF .SR_VALUE = 1'b0;
    defparam \lcd_de~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_dv~FF  (.D(\u_lcd_driver/n133 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_dv )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_dv~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_dv~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[0]~FF  (.D(\u_lcd_driver/n34 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[1]~FF  (.D(\u_lcd_driver/n82 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[2]~FF  (.D(\u_lcd_driver/n81 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[3]~FF  (.D(\u_lcd_driver/n80 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[4]~FF  (.D(\u_lcd_driver/n79 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[5]~FF  (.D(\u_lcd_driver/n78 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[6]~FF  (.D(\u_lcd_driver/n77 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[7]~FF  (.D(\u_lcd_driver/n76 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[8]~FF  (.D(\u_lcd_driver/n75 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[9]~FF  (.D(\u_lcd_driver/n74 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[10]~FF  (.D(\u_lcd_driver/n73 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[11]~FF  (.D(\u_lcd_driver/n72 ), .CE(\u_lcd_driver/equal_17/n23 ), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/vcnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(108)
    defparam \u_lcd_driver/vcnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22  (.D(n7351), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13  (.D(n7326), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[5]~FF  (.D(\lcd_data[5] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[1]~FF  (.D(\u_lcd_driver/n33 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[2]~FF  (.D(\u_lcd_driver/n32 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[3]~FF  (.D(\u_lcd_driver/n31 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[4]~FF  (.D(\u_lcd_driver/n30 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[5]~FF  (.D(\u_lcd_driver/n29 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[6]~FF  (.D(\u_lcd_driver/n28 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[7]~FF  (.D(\u_lcd_driver/n27 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[8]~FF  (.D(\u_lcd_driver/n26 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[9]~FF  (.D(\u_lcd_driver/n25 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[10]~FF  (.D(\u_lcd_driver/n24 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[11]~FF  (.D(\u_lcd_driver/n23 ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(r_hdmi_rst_n), .Q(\u_lcd_driver/hcnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(87)
    defparam \u_lcd_driver/hcnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[0]~FF  (.D(\u_rgb2dvi/enc_0/n869 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[0]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[0]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[0]~FF  (.D(n3195), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_0/acc[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[1]~FF  (.D(\u_rgb2dvi/enc_0/n764 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[1]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[1]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[1]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[1]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[1]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[1]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[2]~FF  (.D(\u_rgb2dvi/enc_0/n770 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[2]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[2]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[2]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[2]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[2]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[3]~FF  (.D(\u_rgb2dvi/enc_0/n776 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[3]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[3]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[3]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[3]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[3]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[3]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[4]~FF  (.D(\u_rgb2dvi/enc_0/n782 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[4]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[4]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[4]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[5]~FF  (.D(\u_rgb2dvi/enc_0/n788 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[5]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[5]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[5]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[5]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[5]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[5]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[6]~FF  (.D(\u_rgb2dvi/enc_0/n794 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[6]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[6]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[6]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[6]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[6]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[6]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[7]~FF  (.D(\u_rgb2dvi/enc_0/n800 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[7]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[7]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[7]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[7]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[7]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[7]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[8]~FF  (.D(\u_rgb2dvi/enc_0/n806 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[8]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[8]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[8]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd0[9]~FF  (.D(\u_rgb2dvi/enc_0/n812 ), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\w_hdmi_txd0[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd0[9]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .SR_POLARITY = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd0[9]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd0[9]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd0[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[1]~FF  (.D(n376), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_0/acc[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[2]~FF  (.D(n374), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_0/acc[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[3]~FF  (.D(n372), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_0/acc[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_0/acc[4]~FF  (.D(n371), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_0/acc[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_0/acc[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[0]~FF  (.D(\u_rgb2dvi/enc_1/q_out[0] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[0]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[0]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[0]~FF  (.D(n3254), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_1/acc[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[1]~FF  (.D(\u_rgb2dvi/enc_1/q_out[1] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[1]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[1]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[1]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[1]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[1]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[2]~FF  (.D(\u_rgb2dvi/enc_1/q_out[2] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[2]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[2]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[2]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[2]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[2]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[3]~FF  (.D(\u_rgb2dvi/enc_1/q_out[3] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[3]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[3]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[3]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[3]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[3]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[4]~FF  (.D(\u_rgb2dvi/enc_1/q_out[4] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[4]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[4]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[4]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[4]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[4]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[5]~FF  (.D(\u_rgb2dvi/enc_1/q_out[5] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[5]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[5]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[5]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[5]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[5]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[6]~FF  (.D(\u_rgb2dvi/enc_1/q_out[6] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[6]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[6]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[6]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[6]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[6]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[7]~FF  (.D(\u_rgb2dvi/enc_1/q_out[7] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[7]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[7]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[7]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[7]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[7]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[8]~FF  (.D(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[8]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[8]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd1[9]~FF  (.D(\u_rgb2dvi/enc_1/q_out[9] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[9]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd1[9]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[9]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd1[9]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd1[9]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[1]~FF  (.D(n350), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_1/acc[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[2]~FF  (.D(n348), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_1/acc[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[3]~FF  (.D(n346), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_1/acc[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_1/acc[4]~FF  (.D(n345), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_1/acc[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_1/acc[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[0]~FF  (.D(\u_rgb2dvi/enc_2/q_out[0] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[0]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[0]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[0]~FF  (.D(n3331), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_2/acc[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[1]~FF  (.D(\u_rgb2dvi/enc_2/q_out[1] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[1]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[1]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[1]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[1]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[1]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[2]~FF  (.D(\u_rgb2dvi/enc_2/q_out[2] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[2]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[2]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[2]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[2]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[2]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[3]~FF  (.D(\u_rgb2dvi/enc_2/q_out[3] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[3]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[3]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[3]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[3]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[3]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[4]~FF  (.D(\u_rgb2dvi/enc_2/q_out[4] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[4]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[4]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[4]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[4]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[4]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[5]~FF  (.D(\u_rgb2dvi/enc_2/q_out[5] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[5]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[5]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[5]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[5]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[5]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[6]~FF  (.D(\u_rgb2dvi/enc_2/q_out[6] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[6]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[6]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[6]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[6]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[6]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[7]~FF  (.D(\u_rgb2dvi/enc_2/q_out[7] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[7]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[7]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[7]~FF .D_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[7]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[7]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \w_hdmi_txd2[9]~FF  (.D(\u_rgb2dvi/enc_2/q_out[9] ), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(lcd_de), .Q(\w_hdmi_txd2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(167)
    defparam \w_hdmi_txd2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[9]~FF .CE_POLARITY = 1'b1;
    defparam \w_hdmi_txd2[9]~FF .SR_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[9]~FF .D_POLARITY = 1'b0;
    defparam \w_hdmi_txd2[9]~FF .SR_SYNC = 1'b1;
    defparam \w_hdmi_txd2[9]~FF .SR_VALUE = 1'b0;
    defparam \w_hdmi_txd2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[1]~FF  (.D(n341), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_2/acc[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[2]~FF  (.D(n339), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_2/acc[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[3]~FF  (.D(n337), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_2/acc[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_rgb2dvi/enc_2/acc[4]~FF  (.D(n336), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(lcd_de), .Q(\u_rgb2dvi/enc_2/acc[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .D_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_SYNC = 1'b1;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_VALUE = 1'b0;
    defparam \u_rgb2dvi/enc_2/acc[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_txc_o[1]~FF  (.D(\r_hdmi_txc_o[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(hdmi_txc_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_txc_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_txc_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_txc_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_txc_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_txc_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_txc_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_txc_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_txc_o[9]~FF  (.D(rc_hdmi_tx), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(\r_hdmi_txc_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_txc_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .SR_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_txc_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_txc_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[1]~FF  (.D(n591), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx0_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[2]~FF  (.D(n590), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx0_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[2]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[3]~FF  (.D(n589), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx0_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[3]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx0_o[4]~FF  (.D(n588), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx0_o[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx0_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx0_o[4]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx0_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[5]~FF  (.D(\w_hdmi_txd0[5] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx0_o[5]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[5]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[5]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[5]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[5]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[5]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[6]~FF  (.D(\w_hdmi_txd0[6] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx0_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[6]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[6]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[6]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[7]~FF  (.D(\w_hdmi_txd0[7] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx0_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[7]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[7]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[8]~FF  (.D(\w_hdmi_txd0[8] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx0_o[8]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[8]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[8]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[8]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[8]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[8]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx0_o[9]~FF  (.D(\w_hdmi_txd0[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx0_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx0_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx0_o[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[9]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx0_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx0_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx0_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[1]~FF  (.D(n602_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx1_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[2]~FF  (.D(n601_2), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx1_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[2]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[3]~FF  (.D(n600), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx1_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[3]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx1_o[4]~FF  (.D(n599), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx1_o[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx1_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx1_o[4]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx1_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[5]~FF  (.D(\w_hdmi_txd1[5] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx1_o[5]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[5]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[5]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[5]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[5]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[5]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[6]~FF  (.D(\w_hdmi_txd1[6] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx1_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[6]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[6]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[6]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[7]~FF  (.D(\w_hdmi_txd1[7] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx1_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[7]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[7]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[8]~FF  (.D(\w_hdmi_txd1[8] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx1_o[8]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[8]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[8]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[8]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[8]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[8]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx1_o[9]~FF  (.D(\w_hdmi_txd1[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx1_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx1_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx1_o[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[9]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx1_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx1_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx1_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[1]~FF  (.D(n613), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx2_o[1]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[1]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[2]~FF  (.D(n612), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx2_o[2]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[2]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[3]~FF  (.D(n611), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx2_o[3]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[3]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hdmi_tx2_o[4]~FF  (.D(n610), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(1'b0), .Q(hdmi_tx2_o[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \hdmi_tx2_o[4]~FF .CLK_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .CE_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .SR_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .D_POLARITY = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .SR_SYNC = 1'b1;
    defparam \hdmi_tx2_o[4]~FF .SR_VALUE = 1'b0;
    defparam \hdmi_tx2_o[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[5]~FF  (.D(\w_hdmi_txd2[5] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx2_o[5]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[5]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[5]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[5]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[5]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[5]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[6]~FF  (.D(\w_hdmi_txd2[6] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx2_o[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[6]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[6]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[6]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[7]~FF  (.D(\w_hdmi_txd2[7] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx2_o[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[7]~FF .D_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[7]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_hdmi_tx2_o[9]~FF  (.D(\w_hdmi_txd2[9] ), .CE(1'b1), .CLK(\hdmi_clk2x_i~O ), 
           .SR(rc_hdmi_tx), .Q(\r_hdmi_tx2_o[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(545)
    defparam \r_hdmi_tx2_o[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_hdmi_tx2_o[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[9]~FF .D_POLARITY = 1'b0;
    defparam \r_hdmi_tx2_o[9]~FF .SR_SYNC = 1'b1;
    defparam \r_hdmi_tx2_o[9]~FF .SR_VALUE = 1'b0;
    defparam \r_hdmi_tx2_o[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[1]~FF  (.D(n3471), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[2]~FF  (.D(n3469), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[3]~FF  (.D(n3467), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[4]~FF  (.D(n3465), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[5]~FF  (.D(n3429), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[6]~FF  (.D(n3427), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[7]~FF  (.D(n3426), .CE(n9_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(121)
    defparam \PowerOnResetCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] ), 
            .I1(1'b0), .CI(n7562), .O(n176), .CO(n177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i2  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0] ), .CI(1'b0), 
            .O(n197), .CO(n198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i2 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i2  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] ), .CI(1'b0), 
            .O(n219), .CO(n220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i2 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i2  (.I0(\i2c_config_index[1] ), 
            .I1(\i2c_config_index[0] ), .CI(1'b0), .O(n222), .CO(n223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i2 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i5  (.I0(\u_rgb2dvi/enc_2/acc[4] ), .I1(n3881), 
            .CI(n338), .O(n336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i4  (.I0(\u_rgb2dvi/enc_2/acc[3] ), .I1(n3884), 
            .CI(n340), .O(n337), .CO(n338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i3  (.I0(\u_rgb2dvi/enc_2/acc[2] ), .I1(n3887), 
            .CI(n342), .O(n339), .CO(n340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i2  (.I0(\u_rgb2dvi/enc_2/acc[1] ), .I1(n3890), 
            .CI(n3332), .O(n341), .CO(n342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_75/i4  (.I0(n358), .I1(1'b0), .CI(n380), 
            .O(n343), .CO(n344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_2/add_75/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_75/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i5  (.I0(\u_rgb2dvi/enc_1/acc[4] ), .I1(n3895), 
            .CI(n347), .O(n345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i4  (.I0(\u_rgb2dvi/enc_1/acc[3] ), .I1(n3898), 
            .CI(n349), .O(n346), .CO(n347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i3  (.I0(\u_rgb2dvi/enc_1/acc[2] ), .I1(n3901), 
            .CI(n351), .O(n348), .CO(n349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i2  (.I0(\u_rgb2dvi/enc_1/acc[1] ), .I1(n3904), 
            .CI(n3255), .O(n350), .CO(n351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i5  (.I0(n364), .I1(1'b1), .CI(n354), 
            .O(n352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i4  (.I0(n365), .I1(1'b1), .CI(n356), 
            .O(n353), .CO(n354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i3  (.I0(n367), .I1(1'b1), .CI(n3208), 
            .O(n355), .CO(n356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i5  (.I0(1'b0), .I1(1'b1), .CI(n359), 
            .O(n357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i4  (.I0(n3913), .I1(n3923), .CI(n361), 
            .O(n358), .CO(n359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i3  (.I0(n3916), .I1(n3926), .CI(n363), 
            .O(n360), .CO(n361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/sub_52/add_2/i2  (.I0(n3919), .I1(n3920), .CI(n7579), 
            .O(n362), .CO(n363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(79)
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_52/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i5  (.I0(1'b0), .I1(1'b1), .CI(n366), 
            .O(n364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i4  (.I0(n3923), .I1(n3913), .CI(n368), 
            .O(n365), .CO(n366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i3  (.I0(n3926), .I1(n3916), .CI(n370), 
            .O(n367), .CO(n368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/sub_50/add_2/i2  (.I0(n3920), .I1(n3919), .CI(n7578), 
            .O(n369), .CO(n370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i2 .I0_POLARITY = 1'b0;
    defparam \u_rgb2dvi/enc_0/sub_50/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i5  (.I0(\u_rgb2dvi/enc_0/acc[4] ), .I1(n3932), 
            .CI(n373), .O(n371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i4  (.I0(\u_rgb2dvi/enc_0/acc[3] ), .I1(n3935), 
            .CI(n375), .O(n372), .CO(n373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i3  (.I0(\u_rgb2dvi/enc_0/acc[2] ), .I1(n3938), 
            .CI(n377), .O(n374), .CO(n375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i2  (.I0(\u_rgb2dvi/enc_0/acc[1] ), .I1(n3941), 
            .CI(n3196), .O(n376), .CO(n377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_75/i5  (.I0(n357), .I1(1'b0), .CI(n344), 
            .O(n378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_0/add_75/i5 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_75/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_75/i3  (.I0(n360), .I1(1'b0), .CI(n3040), 
            .O(n379), .CO(n380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_0/add_75/i3 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_75/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i12  (.I0(\u_lcd_driver/vcnt[11] ), .I1(1'b0), 
            .CI(n383), .O(n381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i12 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i11  (.I0(\u_lcd_driver/vcnt[10] ), .I1(1'b0), 
            .CI(n385), .O(n382), .CO(n383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i11 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i10  (.I0(\u_lcd_driver/vcnt[9] ), .I1(1'b0), 
            .CI(n387), .O(n384), .CO(n385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i10 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i9  (.I0(\u_lcd_driver/vcnt[8] ), .I1(1'b0), 
            .CI(n389), .O(n386), .CO(n387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i9 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i8  (.I0(\u_lcd_driver/vcnt[7] ), .I1(1'b0), 
            .CI(n391), .O(n388), .CO(n389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i8 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i7  (.I0(\u_lcd_driver/vcnt[6] ), .I1(1'b0), 
            .CI(n393), .O(n390), .CO(n391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i7 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i6  (.I0(\u_lcd_driver/vcnt[5] ), .I1(1'b0), 
            .CI(n395), .O(n392), .CO(n393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i6 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i5  (.I0(\u_lcd_driver/vcnt[4] ), .I1(1'b0), 
            .CI(n397), .O(n394), .CO(n395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i5 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i4  (.I0(\u_lcd_driver/vcnt[3] ), .I1(1'b0), 
            .CI(n399), .O(n396), .CO(n397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i4 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i3  (.I0(\u_lcd_driver/vcnt[2] ), .I1(1'b0), 
            .CI(n3030), .O(n398), .CO(n399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i3 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i12  (.I0(\u_lcd_driver/hcnt[11] ), .I1(1'b0), 
            .CI(n402), .O(n400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i12 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i11  (.I0(\u_lcd_driver/hcnt[10] ), .I1(1'b0), 
            .CI(n404), .O(n401), .CO(n402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i11 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i10  (.I0(\u_lcd_driver/hcnt[9] ), .I1(1'b0), 
            .CI(n406), .O(n403), .CO(n404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i10 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i9  (.I0(\u_lcd_driver/hcnt[8] ), .I1(1'b0), 
            .CI(n408), .O(n405), .CO(n406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i9 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i8  (.I0(\u_lcd_driver/hcnt[7] ), .I1(1'b0), 
            .CI(n410), .O(n407), .CO(n408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i8 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i7  (.I0(\u_lcd_driver/hcnt[6] ), .I1(1'b0), 
            .CI(n412), .O(n409), .CO(n410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i7 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i6  (.I0(\u_lcd_driver/hcnt[5] ), .I1(1'b0), 
            .CI(n414), .O(n411), .CO(n412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i6 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i5  (.I0(\u_lcd_driver/hcnt[4] ), .I1(1'b0), 
            .CI(n416), .O(n413), .CO(n414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i5 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i4  (.I0(\u_lcd_driver/hcnt[3] ), .I1(1'b0), 
            .CI(n418), .O(n415), .CO(n416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i4 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i3  (.I0(\u_lcd_driver/hcnt[2] ), .I1(1'b0), 
            .CI(n2538), .O(n417), .CO(n418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i3 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i8  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] ), 
            .CI(n421), .O(n419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i7  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] ), 
            .CI(n423), .O(n420), .CO(n421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i6  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] ), 
            .CI(n425), .O(n422), .CO(n423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i5  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .CI(n427), .O(n424), .CO(n425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i4  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .CI(n429), .O(n426), .CO(n427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i3  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .CI(n431), .O(n428), .CO(n429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i2  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .CI(n2521), .O(n430), .CO(n431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i2  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[1] ), 
            .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[0] ), .CI(1'b0), .O(n443), 
            .CO(n444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i2 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i13  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] ), 
            .I1(1'b0), .CI(n465), .O(n457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i12  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] ), 
            .I1(1'b0), .CI(n467), .O(n464), .CO(n465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i11  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), 
            .I1(1'b0), .CI(n480), .O(n466), .CO(n467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i10  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), 
            .I1(1'b0), .CI(n525), .O(n479), .CO(n480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i9  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
            .I1(1'b0), .CI(n535), .O(n524), .CO(n525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i8  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I1(1'b0), .CI(n537), .O(n534), .CO(n535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i7  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I1(1'b0), .CI(n539), .O(n536), .CO(n537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i6  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I1(1'b0), .CI(n541), .O(n538), .CO(n539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i5  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I1(1'b0), .CI(n543), .O(n540), .CO(n541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i4  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] ), 
            .I1(1'b0), .CI(n545), .O(n542), .CO(n543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i3  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] ), 
            .I1(1'b0), .CI(n2518), .O(n544), .CO(n545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i9  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I1(1'b0), .CI(n548), .O(n546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i8  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(1'b0), .CI(n550), .O(n547), .CO(n548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i7  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(1'b0), .CI(n552), .O(n549), .CO(n550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i6  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(1'b0), .CI(n554), .O(n551), .CO(n552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i5  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(1'b0), .CI(n556), .O(n553), .CO(n554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i4  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(1'b0), .CI(n2511), .O(n555), .CO(n556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] ), 
            .I1(n4132), .CI(n559), .O(n557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] ), 
            .I1(n4135), .CI(n561), .O(n558), .CO(n559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] ), 
            .I1(n4138), .CI(n597), .CO(n561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i2  (.I0(\u_sensor_frame_count/delay_cnt[1] ), 
            .I1(\u_sensor_frame_count/delay_cnt[0] ), .CI(1'b0), .O(n575), 
            .CO(n576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i2 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .I1(n4176), .CI(n629), .CO(n597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i2  (.I0(\u_sensor_frame_count/cmos_fps_cnt[1] ), 
            .I1(\u_sensor_frame_count/cmos_fps_cnt[0] ), .CI(1'b0), .O(n601), 
            .CO(n602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i2 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i4  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .I1(n4211), .CI(n639), .CO(n629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i3  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .I1(n4222), .CI(n641), .CO(n639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i2  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I1(n4225), .CI(n2367), .CO(n641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14  (.I0(1'b0), 
            .I1(1'b1), .CI(n644), .O(n642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .CI(n646), .O(n643), .CO(n644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), .CI(n648), 
            .O(n645), .CO(n646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), .CI(n650), 
            .O(n647), .CO(n648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), .CI(n652), 
            .O(n649), .CO(n650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), .CI(n654), 
            .O(n651), .CO(n652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), .CI(n656), 
            .O(n653), .CO(n654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), .CI(n658), 
            .O(n655), .CO(n656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), .CI(n2356), 
            .O(n657), .CO(n658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I1(1'b0), .CI(n661), .O(n659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I1(1'b0), .CI(n663), .O(n660), .CO(n661)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I1(1'b0), .CI(n665), .O(n662), .CO(n663)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I1(1'b0), .CI(n667), .O(n664), .CO(n665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I1(1'b0), .CI(n669), .O(n666), .CO(n667)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), 
            .I1(1'b0), .CI(n671), .O(n668), .CO(n669)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), 
            .I1(1'b0), .CI(n2350), .O(n670), .CO(n671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
            .I1(1'b0), .CI(n684), .O(n672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/waddr[0] ), .CI(1'b0), .O(n681), 
            .CO(n682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), 
            .I1(1'b0), .CI(n713), .O(n683), .CO(n684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[2] ), 
            .I1(1'b0), .CI(n682), .O(n703), .CO(n704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), 
            .I1(1'b0), .CI(n719), .O(n712), .CO(n713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[0] ), .CI(1'b0), .O(n715), 
            .CO(n716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), 
            .I1(1'b0), .CI(n724), .O(n718), .CO(n719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1  (.I0(n4296), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[0] ), .CI(n7563), .O(n721), 
            .CO(n722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), 
            .I1(1'b0), .CI(n738), .O(n723), .CO(n724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i2  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0] ), .CI(1'b0), 
            .O(n735), .CO(n736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(1'b0), .CI(n740), .O(n737), .CO(n738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(1'b0), .CI(n742), .O(n739), .CO(n740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(1'b0), .CI(n744), .O(n741), .CO(n742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(1'b0), .CI(n746), .O(n743), .CO(n744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(1'b0), .CI(n2270), .O(n745), .CO(n746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i14  (.I0(\u_axi4_ctrl/araddr[23] ), .I1(1'b0), 
            .CI(n749), .O(n747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i14 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i13  (.I0(\u_axi4_ctrl/araddr[22] ), .I1(1'b0), 
            .CI(n751), .O(n748), .CO(n749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i12  (.I0(\u_axi4_ctrl/araddr[21] ), .I1(1'b0), 
            .CI(n753), .O(n750), .CO(n751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i11  (.I0(\u_axi4_ctrl/araddr[20] ), .I1(1'b0), 
            .CI(n755), .O(n752), .CO(n753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i10  (.I0(\u_axi4_ctrl/araddr[19] ), .I1(1'b0), 
            .CI(n770), .O(n754), .CO(n755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i9  (.I0(\u_axi4_ctrl/araddr[18] ), .I1(1'b0), 
            .CI(n772), .O(n769), .CO(n770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i8  (.I0(\u_axi4_ctrl/araddr[17] ), .I1(1'b0), 
            .CI(n774), .O(n771), .CO(n772)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i7  (.I0(\u_axi4_ctrl/araddr[16] ), .I1(1'b0), 
            .CI(n776), .O(n773), .CO(n774)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i6  (.I0(\u_axi4_ctrl/araddr[15] ), .I1(1'b0), 
            .CI(n778), .O(n775), .CO(n776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i5  (.I0(\u_axi4_ctrl/araddr[14] ), .I1(1'b0), 
            .CI(n780), .O(n777), .CO(n778)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i4  (.I0(\u_axi4_ctrl/araddr[13] ), .I1(1'b0), 
            .CI(n2189), .O(n779), .CO(n780)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i14  (.I0(\u_axi4_ctrl/awaddr[23] ), .I1(1'b0), 
            .CI(n783), .O(n781)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i14 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i13  (.I0(\u_axi4_ctrl/awaddr[22] ), .I1(1'b0), 
            .CI(n785), .O(n782), .CO(n783)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i12  (.I0(\u_axi4_ctrl/awaddr[21] ), .I1(1'b0), 
            .CI(n787), .O(n784), .CO(n785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i11  (.I0(\u_axi4_ctrl/awaddr[20] ), .I1(1'b0), 
            .CI(n789), .O(n786), .CO(n787)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i10  (.I0(\u_axi4_ctrl/awaddr[19] ), .I1(1'b0), 
            .CI(n791), .O(n788), .CO(n789)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i9  (.I0(\u_axi4_ctrl/awaddr[18] ), .I1(1'b0), 
            .CI(n793), .O(n790), .CO(n791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i8  (.I0(\u_axi4_ctrl/awaddr[17] ), .I1(1'b0), 
            .CI(n795), .O(n792), .CO(n793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i7  (.I0(\u_axi4_ctrl/awaddr[16] ), .I1(1'b0), 
            .CI(n797), .O(n794), .CO(n795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i6  (.I0(\u_axi4_ctrl/awaddr[15] ), .I1(1'b0), 
            .CI(n799), .O(n796), .CO(n797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i5  (.I0(\u_axi4_ctrl/awaddr[14] ), .I1(1'b0), 
            .CI(n801), .O(n798), .CO(n799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i4  (.I0(\u_axi4_ctrl/awaddr[13] ), .I1(1'b0), 
            .CI(n803), .O(n800), .CO(n801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i3  (.I0(\u_axi4_ctrl/awaddr[12] ), .I1(1'b0), 
            .CI(n2150), .O(n802), .CO(n803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i2  (.I0(\u_scaler_gray/vs_cnt[1] ), .I1(\u_scaler_gray/vs_cnt[0] ), 
            .CI(1'b0), .O(n900), .CO(n901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i2  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] ), .CI(1'b0), 
            .O(n904), .CO(n905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i2  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_addra[0] ), .CI(1'b0), 
            .O(n911), .CO(n912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i2  (.I0(\u_scaler_gray/destx[1] ), 
            .I1(\u_scaler_gray/destx[0] ), .CI(1'b0), .O(n916), .CO(n917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21] ), 
            .I1(1'b0), .CI(n921), .O(n919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20] ), 
            .I1(1'b0), .CI(n923), .O(n920), .CO(n921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19] ), 
            .I1(1'b0), .CI(n925), .O(n922), .CO(n923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18] ), 
            .I1(1'b0), .CI(n927), .O(n924), .CO(n925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17] ), 
            .I1(1'b0), .CI(n931), .O(n926), .CO(n927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16] ), 
            .I1(1'b0), .CI(n933), .O(n930), .CO(n931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15] ), 
            .I1(1'b0), .CI(n937), .O(n932), .CO(n933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i2  (.I0(\u_scaler_gray/desty[1] ), 
            .I1(\u_scaler_gray/desty[0] ), .CI(1'b0), .O(n934), .CO(n935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14] ), 
            .I1(1'b0), .CI(n1914), .O(n936), .CO(n937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[20] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[20] ), 
            .CI(n943), .O(n940), .CO(n7564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[19] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[19] ), 
            .CI(n945), .O(n942), .CO(n943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[18] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[18] ), 
            .CI(n947), .O(n944), .CO(n945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[17] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[17] ), 
            .CI(n949), .O(n946), .CO(n947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[16] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[16] ), 
            .CI(n951), .O(n948), .CO(n949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[15] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[15] ), 
            .CI(n953), .O(n950), .CO(n951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[14] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[14] ), 
            .CI(n955), .O(n952), .CO(n953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[13] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[13] ), 
            .CI(n957), .O(n954), .CO(n955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[12] ), 
            .CI(n959), .O(n956), .CO(n957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[11] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[11] ), 
            .CI(n960), .O(n958), .CO(n959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[10] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[10] ), 
            .CI(n961), .CO(n960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[9] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[9] ), 
            .CI(n962), .CO(n961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[8] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[8] ), 
            .CI(n965), .CO(n962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[7] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[7] ), 
            .CI(n973), .CO(n965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[6] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[6] ), 
            .CI(n974), .CO(n973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[5] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[5] ), 
            .CI(n1008), .CO(n974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[4] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[4] ), 
            .CI(n1009), .CO(n1008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[3] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[3] ), 
            .CI(n1010), .CO(n1009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[2] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[2] ), 
            .CI(n1011), .CO(n1010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[1] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[1] ), 
            .CI(n1910), .CO(n1011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[19] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[19] ), 
            .CI(n1015), .O(n1012), .CO(n7565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[18] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[18] ), 
            .CI(n1017), .O(n1014), .CO(n1015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[17] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[17] ), 
            .CI(n1019), .O(n1016), .CO(n1017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[16] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[16] ), 
            .CI(n1021), .O(n1018), .CO(n1019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[15] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[15] ), 
            .CI(n1023), .O(n1020), .CO(n1021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[14] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[14] ), 
            .CI(n1025), .O(n1022), .CO(n1023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[13] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[13] ), 
            .CI(n1027), .O(n1024), .CO(n1025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[12] ), 
            .CI(n1029), .O(n1026), .CO(n1027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[11] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[11] ), 
            .CI(n1031), .O(n1028), .CO(n1029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[10] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[10] ), 
            .CI(n1033), .O(n1030), .CO(n1031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[9] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[9] ), 
            .CI(n1035), .O(n1032), .CO(n1033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[8] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[8] ), 
            .CI(n1037), .O(n1034), .CO(n1035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[7] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[7] ), 
            .CI(n1039), .O(n1036), .CO(n1037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[6] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[6] ), 
            .CI(n1041), .O(n1038), .CO(n1039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[5] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[5] ), 
            .CI(n1043), .O(n1040), .CO(n1041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[4] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[4] ), 
            .CI(n1045), .O(n1042), .CO(n1043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[3] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[3] ), 
            .CI(n1047), .O(n1044), .CO(n1045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[2] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[2] ), 
            .CI(n1049), .O(n1046), .CO(n1047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[1] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[1] ), 
            .CI(n1909), .O(n1048), .CO(n1049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[19] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[19] ), 
            .CI(n1068), .O(n1065), .CO(n7566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[18] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[18] ), 
            .CI(n1070), .O(n1067), .CO(n1068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[17] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[17] ), 
            .CI(n1072), .O(n1069), .CO(n1070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[16] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[16] ), 
            .CI(n1074), .O(n1071), .CO(n1072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[15] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[15] ), 
            .CI(n1076), .O(n1073), .CO(n1074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[14] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[14] ), 
            .CI(n1078), .O(n1075), .CO(n1076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[13] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[13] ), 
            .CI(n1080), .O(n1077), .CO(n1078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[12] ), 
            .CI(n1082), .O(n1079), .CO(n1080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[11] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[11] ), 
            .CI(n1084), .O(n1081), .CO(n1082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[10] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[10] ), 
            .CI(n1086), .O(n1083), .CO(n1084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[9] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[9] ), 
            .CI(n1088), .O(n1085), .CO(n1086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[8] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[8] ), 
            .CI(n1090), .O(n1087), .CO(n1088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[7] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[7] ), 
            .CI(n1092), .O(n1089), .CO(n1090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[6] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[6] ), 
            .CI(n1094), .O(n1091), .CO(n1092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[5] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[5] ), 
            .CI(n1096), .O(n1093), .CO(n1094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[4] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[4] ), 
            .CI(n1098), .O(n1095), .CO(n1096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[3] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[3] ), 
            .CI(n1100), .O(n1097), .CO(n1098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[2] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[2] ), 
            .CI(n1102), .O(n1099), .CO(n1100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[1] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[1] ), 
            .CI(n1740), .O(n1101), .CO(n1102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[23] ), 
            .I1(1'b0), .CI(n1105), .O(n1103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[22] ), 
            .I1(1'b0), .CI(n1107), .O(n1104), .CO(n1105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[21] ), 
            .I1(1'b0), .CI(n1109), .O(n1106), .CO(n1107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[20] ), 
            .I1(1'b0), .CI(n1111), .O(n1108), .CO(n1109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[19] ), 
            .I1(1'b0), .CI(n1115), .O(n1110), .CO(n1111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[18] ), 
            .I1(1'b0), .CI(n1133), .O(n1114), .CO(n1115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[17] ), 
            .I1(1'b0), .CI(n1135), .O(n1132), .CO(n1133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[16] ), 
            .I1(1'b0), .CI(n1137), .O(n1134), .CO(n1135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[15] ), 
            .I1(1'b0), .CI(n1139), .O(n1136), .CO(n1137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[14] ), 
            .I1(1'b0), .CI(n1141), .O(n1138), .CO(n1139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[13] ), 
            .I1(1'b0), .CI(n1724), .O(n1140), .CO(n1141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[23] ), 
            .I1(1'b0), .CI(n1144), .O(n1142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[22] ), 
            .I1(1'b0), .CI(n1146), .O(n1143), .CO(n1144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[21] ), 
            .I1(1'b0), .CI(n1148), .O(n1145), .CO(n1146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[20] ), 
            .I1(1'b0), .CI(n1150), .O(n1147), .CO(n1148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[19] ), 
            .I1(1'b0), .CI(n1152), .O(n1149), .CO(n1150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[18] ), 
            .I1(1'b0), .CI(n1154), .O(n1151), .CO(n1152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[17] ), 
            .I1(1'b0), .CI(n1156), .O(n1153), .CO(n1154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[16] ), 
            .I1(1'b0), .CI(n1158), .O(n1155), .CO(n1156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[15] ), 
            .I1(1'b0), .CI(n1160), .O(n1157), .CO(n1158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[14] ), 
            .I1(1'b0), .CI(n1162), .O(n1159), .CO(n1160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[13] ), 
            .I1(1'b0), .CI(n1722), .O(n1161), .CO(n1162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[23] ), 
            .I1(1'b0), .CI(n1165), .O(n1163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[22] ), 
            .I1(1'b0), .CI(n1167), .O(n1164), .CO(n1165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[21] ), 
            .I1(1'b0), .CI(n1169), .O(n1166), .CO(n1167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[20] ), 
            .I1(1'b0), .CI(n1171), .O(n1168), .CO(n1169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[19] ), 
            .I1(1'b0), .CI(n1173), .O(n1170), .CO(n1171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[18] ), 
            .I1(1'b0), .CI(n1175), .O(n1172), .CO(n1173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[17] ), 
            .I1(1'b0), .CI(n1177), .O(n1174), .CO(n1175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[16] ), 
            .I1(1'b0), .CI(n1179), .O(n1176), .CO(n1177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[15] ), 
            .I1(1'b0), .CI(n1181), .O(n1178), .CO(n1179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[14] ), 
            .I1(1'b0), .CI(n1183), .O(n1180), .CO(n1181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[13] ), 
            .I1(1'b0), .CI(n1720), .O(n1182), .CO(n1183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[23] ), 
            .I1(1'b0), .CI(n1201), .O(n1199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[22] ), 
            .I1(1'b0), .CI(n1203), .O(n1200), .CO(n1201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[21] ), 
            .I1(1'b0), .CI(n1205), .O(n1202), .CO(n1203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[20] ), 
            .I1(1'b0), .CI(n1207), .O(n1204), .CO(n1205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[19] ), 
            .I1(1'b0), .CI(n1209), .O(n1206), .CO(n1207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[18] ), 
            .I1(1'b0), .CI(n1211), .O(n1208), .CO(n1209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[17] ), 
            .I1(1'b0), .CI(n1213), .O(n1210), .CO(n1211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[16] ), 
            .I1(1'b0), .CI(n1215), .O(n1212), .CO(n1213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[15] ), 
            .I1(1'b0), .CI(n1217), .O(n1214), .CO(n1215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[14] ), 
            .I1(1'b0), .CI(n1219), .O(n1216), .CO(n1217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[13] ), 
            .I1(1'b0), .CI(n1675), .O(n1218), .CO(n1219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i28  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27] ), 
            .I1(1'b1), .CI(n1222), .O(n1220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i27  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26] ), 
            .I1(1'b1), .CI(n1224), .O(n1221), .CO(n1222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i26  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25] ), 
            .I1(1'b1), .CI(n1226), .O(n1223), .CO(n1224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i25  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24] ), 
            .I1(1'b1), .CI(n1228), .O(n1225), .CO(n1226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i24  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23] ), 
            .I1(1'b1), .CI(n1230), .O(n1227), .CO(n1228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i23  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22] ), 
            .I1(1'b1), .CI(n1232), .O(n1229), .CO(n1230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i22  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21] ), 
            .I1(1'b1), .CI(n1234), .O(n1231), .CO(n1232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i21  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20] ), 
            .I1(1'b1), .CI(n1236), .O(n1233), .CO(n1234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19] ), 
            .I1(1'b1), .CI(n1238), .O(n1235), .CO(n1236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18] ), 
            .I1(1'b1), .CI(n1240), .O(n1237), .CO(n1238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17] ), 
            .I1(1'b1), .CI(n1242), .O(n1239), .CO(n1240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16] ), 
            .I1(1'b1), .CI(n1244), .O(n1241), .CO(n1242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15] ), 
            .I1(1'b1), .CI(n1246), .O(n1243), .CO(n1244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14] ), 
            .I1(1'b1), .CI(n1248), .O(n1245), .CO(n1246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13] ), 
            .I1(1'b1), .CI(n1250), .O(n1247), .CO(n1248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12] ), 
            .I1(1'b1), .CI(n1673), .O(n1249), .CO(n1250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i28  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27] ), 
            .CI(n1253), .O(n1251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i27  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26] ), 
            .CI(n1255), .O(n1252), .CO(n1253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i26  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25] ), 
            .CI(n1257), .O(n1254), .CO(n1255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i25  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24] ), 
            .CI(n1259), .O(n1256), .CO(n1257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i24  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23] ), 
            .CI(n1261), .O(n1258), .CO(n1259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i23  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22] ), 
            .CI(n1263), .O(n1260), .CO(n1261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i22  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21] ), 
            .CI(n1265), .O(n1262), .CO(n1263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i21  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20] ), 
            .CI(n1267), .O(n1264), .CO(n1265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i20  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19] ), 
            .CI(n1273), .O(n1266), .CO(n1267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i19  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18] ), 
            .CI(n1275), .O(n1272), .CO(n1273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i18  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17] ), 
            .CI(n1277), .O(n1274), .CO(n1275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i17  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16] ), 
            .CI(n1279), .O(n1276), .CO(n1277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i16  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15] ), 
            .CI(n1281), .O(n1278), .CO(n1279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i15  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14] ), 
            .CI(n1283), .O(n1280), .CO(n1281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i14  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13] ), 
            .CI(n1285), .O(n1282), .CO(n1283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i13  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12] ), 
            .CI(n1287), .O(n1284), .CO(n1285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i12  (.I0(1'b1), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11] ), 
            .CI(n1289), .O(n1286), .CO(n1287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i11  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10] ), 
            .CI(n1291), .O(n1288), .CO(n1289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i10  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9] ), 
            .CI(n1293), .O(n1290), .CO(n1291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i9  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8] ), 
            .CI(n1295), .O(n1292), .CO(n1293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i8  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7] ), 
            .CI(n1297), .O(n1294), .CO(n1295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i7  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6] ), 
            .CI(n1299), .O(n1296), .CO(n1297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i6  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5] ), 
            .CI(n1301), .O(n1298), .CO(n1299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i5  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4] ), 
            .CI(n1303), .O(n1300), .CO(n1301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i4  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3] ), 
            .CI(n1305), .O(n1302), .CO(n1303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i3  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2] ), 
            .CI(n1307), .O(n1304), .CO(n1305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i2  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1] ), 
            .CI(n1643), .O(n1306), .CO(n1307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i28  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27] ), 
            .I1(1'b1), .CI(n1310), .O(n1308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i27  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26] ), 
            .I1(1'b1), .CI(n1312), .O(n1309), .CO(n1310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i26  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25] ), 
            .I1(1'b1), .CI(n1314), .O(n1311), .CO(n1312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i25  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24] ), 
            .I1(1'b1), .CI(n1316), .O(n1313), .CO(n1314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i24  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23] ), 
            .I1(1'b1), .CI(n1318), .O(n1315), .CO(n1316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i23  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22] ), 
            .I1(1'b1), .CI(n1320), .O(n1317), .CO(n1318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i22  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21] ), 
            .I1(1'b1), .CI(n1322), .O(n1319), .CO(n1320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i21  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20] ), 
            .I1(1'b1), .CI(n1324), .O(n1321), .CO(n1322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19] ), 
            .I1(1'b1), .CI(n1326), .O(n1323), .CO(n1324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18] ), 
            .I1(1'b1), .CI(n1328), .O(n1325), .CO(n1326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17] ), 
            .I1(1'b1), .CI(n1352), .O(n1327), .CO(n1328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16] ), 
            .I1(1'b1), .CI(n1354), .O(n1351), .CO(n1352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15] ), 
            .I1(1'b1), .CI(n1356), .O(n1353), .CO(n1354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14] ), 
            .I1(1'b1), .CI(n1358), .O(n1355), .CO(n1356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13] ), 
            .I1(1'b1), .CI(n1360), .O(n1357), .CO(n1358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12] ), 
            .I1(1'b1), .CI(n1641), .O(n1359), .CO(n1360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i28  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27] ), 
            .CI(n1398), .O(n1396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i27  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26] ), 
            .CI(n1400), .O(n1397), .CO(n1398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i26  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25] ), 
            .CI(n1402), .O(n1399), .CO(n1400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i25  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24] ), 
            .CI(n1404), .O(n1401), .CO(n1402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i24  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23] ), 
            .CI(n1406), .O(n1403), .CO(n1404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i23  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22] ), 
            .CI(n1450), .O(n1405), .CO(n1406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i22  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21] ), 
            .CI(n1452), .O(n1449), .CO(n1450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i21  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20] ), 
            .CI(n1454), .O(n1451), .CO(n1452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i21 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i20  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19] ), 
            .CI(n1456), .O(n1453), .CO(n1454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i19  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18] ), 
            .CI(n1458), .O(n1455), .CO(n1456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i18  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17] ), 
            .CI(n1460), .O(n1457), .CO(n1458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i17  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16] ), 
            .CI(n1462), .O(n1459), .CO(n1460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i16  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15] ), 
            .CI(n1464), .O(n1461), .CO(n1462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i15  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14] ), 
            .CI(n1466), .O(n1463), .CO(n1464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i14  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13] ), 
            .CI(n1468), .O(n1465), .CO(n1466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i13  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12] ), 
            .CI(n1470), .O(n1467), .CO(n1468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i12  (.I0(1'b1), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11] ), 
            .CI(n1472), .O(n1469), .CO(n1470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i11  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10] ), 
            .CI(n1474), .O(n1471), .CO(n1472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10  (.I0(1'b0), 
            .I1(DdrCtrl_ALEN_0[0]), .CI(n7567), .O(n1473), .CO(n1474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_15/add_2/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \add_351/i28  (.I0(1'b0), .I1(\u_scaler_gray/destx[15] ), .CI(n1477), 
            .O(n1475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i28 .I0_POLARITY = 1'b1;
    defparam \add_351/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i27  (.I0(1'b0), .I1(\u_scaler_gray/destx[14] ), .CI(n1479), 
            .O(n1476), .CO(n1477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i27 .I0_POLARITY = 1'b1;
    defparam \add_351/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i26  (.I0(\u_scaler_gray/destx[15] ), .I1(\u_scaler_gray/destx[13] ), 
            .CI(n1481), .O(n1478), .CO(n1479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i26 .I0_POLARITY = 1'b1;
    defparam \add_351/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i25  (.I0(\u_scaler_gray/destx[14] ), .I1(\u_scaler_gray/destx[12] ), 
            .CI(n1496), .O(n1480), .CO(n1481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i25 .I0_POLARITY = 1'b1;
    defparam \add_351/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i24  (.I0(\u_scaler_gray/destx[13] ), .I1(\u_scaler_gray/destx[11] ), 
            .CI(n1498), .O(n1495), .CO(n1496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i24 .I0_POLARITY = 1'b1;
    defparam \add_351/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i23  (.I0(\u_scaler_gray/destx[12] ), .I1(\u_scaler_gray/destx[10] ), 
            .CI(n1500), .O(n1497), .CO(n1498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i23 .I0_POLARITY = 1'b1;
    defparam \add_351/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i22  (.I0(\u_scaler_gray/destx[11] ), .I1(\u_scaler_gray/destx[9] ), 
            .CI(n1502), .O(n1499), .CO(n1500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i22 .I0_POLARITY = 1'b1;
    defparam \add_351/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i21  (.I0(\u_scaler_gray/destx[10] ), .I1(\u_scaler_gray/destx[8] ), 
            .CI(n1504), .O(n1501), .CO(n1502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i21 .I0_POLARITY = 1'b1;
    defparam \add_351/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i20  (.I0(\u_scaler_gray/destx[9] ), .I1(\u_scaler_gray/destx[7] ), 
            .CI(n1506), .O(n1503), .CO(n1504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i20 .I0_POLARITY = 1'b1;
    defparam \add_351/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i19  (.I0(\u_scaler_gray/destx[8] ), .I1(\u_scaler_gray/destx[6] ), 
            .CI(n1508), .O(n1505), .CO(n1506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i19 .I0_POLARITY = 1'b1;
    defparam \add_351/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i18  (.I0(\u_scaler_gray/destx[7] ), .I1(\u_scaler_gray/destx[5] ), 
            .CI(n1510), .O(n1507), .CO(n1508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i18 .I0_POLARITY = 1'b1;
    defparam \add_351/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i17  (.I0(\u_scaler_gray/destx[6] ), .I1(\u_scaler_gray/destx[4] ), 
            .CI(n1512), .O(n1509), .CO(n1510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i17 .I0_POLARITY = 1'b1;
    defparam \add_351/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i16  (.I0(\u_scaler_gray/destx[5] ), .I1(\u_scaler_gray/destx[3] ), 
            .CI(n1514), .O(n1511), .CO(n1512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i16 .I0_POLARITY = 1'b1;
    defparam \add_351/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i15  (.I0(\u_scaler_gray/destx[4] ), .I1(\u_scaler_gray/destx[2] ), 
            .CI(n1516), .O(n1513), .CO(n1514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i15 .I0_POLARITY = 1'b1;
    defparam \add_351/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i14  (.I0(\u_scaler_gray/destx[3] ), .I1(\u_scaler_gray/destx[1] ), 
            .CI(n1537), .O(n1515), .CO(n1516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i14 .I0_POLARITY = 1'b1;
    defparam \add_351/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[1] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[0] ), 
            .CI(1'b0), .O(n1534), .CO(n1535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_351/i13  (.I0(\u_scaler_gray/destx[2] ), .I1(\u_scaler_gray/destx[0] ), 
            .CI(1'b0), .O(n1536), .CO(n1537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(54)
    defparam \add_351/i13 .I0_POLARITY = 1'b1;
    defparam \add_351/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11] ), 
            .I1(1'b0), .CI(n7568), .O(n1640), .CO(n1641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(70)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_16/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1  (.I0(1'b0), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0] ), 
            .CI(n7569), .O(n1642), .CO(n1643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(77)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_21/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i28  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[27] ), 
            .I1(1'b0), .CI(n1677), .O(n1671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11] ), 
            .I1(1'b0), .CI(n7570), .O(n1672), .CO(n1673)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(79)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/sub_22/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[11] ), 
            .CI(1'b0), .O(n1674), .CO(n1675)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(65)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_24/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i27  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[26] ), 
            .I1(1'b0), .CI(n1679), .O(n1676), .CO(n1677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i26  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[25] ), 
            .I1(1'b0), .CI(n1681), .O(n1678), .CO(n1679)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i25  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[24] ), 
            .I1(1'b0), .CI(n1683), .O(n1680), .CO(n1681)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i24  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[23] ), 
            .I1(1'b0), .CI(n1685), .O(n1682), .CO(n1683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i23  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[22] ), 
            .I1(1'b0), .CI(n1687), .O(n1684), .CO(n1685)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i22  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[21] ), 
            .I1(1'b0), .CI(n1689), .O(n1686), .CO(n1687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i21  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[20] ), 
            .I1(1'b0), .CI(n1691), .O(n1688), .CO(n1689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[19] ), 
            .I1(1'b0), .CI(n1693), .O(n1690), .CO(n1691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[18] ), 
            .I1(1'b0), .CI(n1714), .O(n1692), .CO(n1693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[17] ), 
            .I1(1'b0), .CI(n1770), .O(n1713), .CO(n1714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[11] ), 
            .CI(1'b0), .O(n1719), .CO(n1720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(66)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_25/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[11] ), 
            .CI(1'b0), .O(n1721), .CO(n1722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(67)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_26/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[11] ), 
            .CI(1'b0), .O(n1723), .CO(n1724)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(68)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/add_27/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[0] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[0] ), 
            .CI(1'b0), .O(n1739), .CO(n1740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(41)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_13/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[16] ), 
            .I1(1'b0), .CI(n2055), .O(n1769), .CO(n1770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[0] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[0] ), 
            .CI(1'b0), .O(n1908), .CO(n1909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(42)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_14/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i1  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add0[0] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level1_add1[0] ), 
            .CI(1'b0), .CO(n1910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(47)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i1 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_18/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i2  (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12] ), 
            .CI(1'b0), .O(n1913), .CO(n1914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(56)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i2 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/add_22/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[15] ), 
            .I1(1'b0), .CI(n2057), .O(n2054), .CO(n2055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[14] ), 
            .I1(1'b0), .CI(n2059), .O(n2056), .CO(n2057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[13] ), 
            .I1(1'b0), .CI(n2061), .O(n2058), .CO(n2059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[12] ), 
            .I1(1'b0), .CI(n2063), .O(n2060), .CO(n2061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[11] ), 
            .I1(1'b1), .CI(n2065), .O(n2062), .CO(n2063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i11  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[10] ), 
            .I1(1'b0), .CI(n2067), .O(n2064), .CO(n2065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i10  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[9] ), 
            .I1(1'b0), .CI(n2108), .O(n2066), .CO(n2067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i9  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[8] ), 
            .I1(1'b1), .CI(n2110), .O(n2107), .CO(n2108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i8  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[7] ), 
            .I1(1'b1), .CI(n2113), .O(n2109), .CO(n2110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i7  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[6] ), 
            .I1(1'b0), .CI(n2116), .O(n2112), .CO(n2113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i6  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[5] ), 
            .I1(1'b0), .CI(n2120), .O(n2115), .CO(n2116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i5  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[4] ), 
            .I1(1'b1), .CI(n2123), .O(n2119), .CO(n2120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i4  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[3] ), 
            .I1(1'b1), .CI(n2127), .O(n2122), .CO(n2123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i2  (.I0(\u_axi4_ctrl/araddr[11] ), .I1(\u_axi4_ctrl/araddr[10] ), 
            .CI(1'b0), .O(n2124), .CO(n2125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i3  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[2] ), 
            .I1(1'b0), .CI(n1535), .O(n2126), .CO(n2127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(62)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i28  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[27] ), 
            .I1(1'b0), .CI(n2134), .O(n2132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i28 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i27  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[26] ), 
            .I1(1'b0), .CI(n2137), .O(n2133), .CO(n2134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i27 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i26  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[25] ), 
            .I1(1'b0), .CI(n2139), .O(n2136), .CO(n2137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i26 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i25  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[24] ), 
            .I1(1'b0), .CI(n2141), .O(n2138), .CO(n2139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i25 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i24  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[23] ), 
            .I1(1'b0), .CI(n2143), .O(n2140), .CO(n2141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i24 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i23  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[22] ), 
            .I1(1'b0), .CI(n2145), .O(n2142), .CO(n2143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i23 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i22  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[21] ), 
            .I1(1'b0), .CI(n2148), .O(n2144), .CO(n2145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i22 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i21  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[20] ), 
            .I1(1'b0), .CI(n2152), .O(n2147), .CO(n2148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i21 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_105/i2  (.I0(\u_axi4_ctrl/awaddr[11] ), .I1(\u_axi4_ctrl/awaddr[10] ), 
            .CI(1'b0), .O(n2149), .CO(n2150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(297)
    defparam \u_axi4_ctrl/add_105/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_105/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i20  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[19] ), 
            .I1(1'b0), .CI(n2154), .O(n2151), .CO(n2152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i20 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i19  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[18] ), 
            .I1(1'b0), .CI(n2156), .O(n2153), .CO(n2154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i19 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i18  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[17] ), 
            .I1(1'b0), .CI(n2159), .O(n2155), .CO(n2156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i18 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i17  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[16] ), 
            .I1(1'b0), .CI(n2161), .O(n2158), .CO(n2159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i17 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i16  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[15] ), 
            .I1(1'b0), .CI(n2163), .O(n2160), .CO(n2161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i15  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[14] ), 
            .I1(1'b0), .CI(n2165), .O(n2162), .CO(n2163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i14  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[13] ), 
            .I1(1'b0), .CI(n2167), .O(n2164), .CO(n2165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i13  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[12] ), 
            .I1(1'b0), .CI(n2170), .O(n2166), .CO(n2167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i12  (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcx_location[11] ), 
            .I1(1'b1), .CI(1'b0), .O(n2169), .CO(n2170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(61)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/add_9/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i16  (.I0(\u_scaler_gray/desty[15] ), 
            .I1(1'b0), .CI(n2225), .O(n2187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_131/i3  (.I0(\u_axi4_ctrl/araddr[12] ), .I1(1'b0), 
            .CI(n2125), .O(n2188), .CO(n2189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/add_131/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_131/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i15  (.I0(\u_scaler_gray/desty[14] ), 
            .I1(1'b0), .CI(n2227), .O(n2224), .CO(n2225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i14  (.I0(\u_scaler_gray/desty[13] ), 
            .I1(1'b0), .CI(n2229), .O(n2226), .CO(n2227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i13  (.I0(\u_scaler_gray/desty[12] ), 
            .I1(1'b0), .CI(n2231), .O(n2228), .CO(n2229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i12  (.I0(\u_scaler_gray/desty[11] ), 
            .I1(1'b0), .CI(n2233), .O(n2230), .CO(n2231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i11  (.I0(\u_scaler_gray/desty[10] ), 
            .I1(1'b0), .CI(n2235), .O(n2232), .CO(n2233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i10  (.I0(\u_scaler_gray/desty[9] ), 
            .I1(1'b0), .CI(n2292), .O(n2234), .CO(n2235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(1'b0), .CI(n2272), .O(n2269), .CO(n2270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] ), .CI(1'b0), 
            .O(n2271), .CO(n2272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i9  (.I0(\u_scaler_gray/desty[8] ), 
            .I1(1'b0), .CI(n2297), .O(n2291), .CO(n2292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i8  (.I0(\u_scaler_gray/desty[7] ), 
            .I1(1'b0), .CI(n2299), .O(n2296), .CO(n2297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i7  (.I0(\u_scaler_gray/desty[6] ), 
            .I1(1'b0), .CI(n2301), .O(n2298), .CO(n2299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i6  (.I0(\u_scaler_gray/desty[5] ), 
            .I1(1'b0), .CI(n2303), .O(n2300), .CO(n2301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i5  (.I0(\u_scaler_gray/desty[4] ), 
            .I1(1'b0), .CI(n2305), .O(n2302), .CO(n2303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i4  (.I0(\u_scaler_gray/desty[3] ), 
            .I1(1'b0), .CI(n2313), .O(n2304), .CO(n2305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_77/i3  (.I0(\u_scaler_gray/desty[2] ), 
            .I1(1'b0), .CI(n935), .O(n2312), .CO(n2313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(209)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_77/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i16  (.I0(\u_scaler_gray/destx[15] ), 
            .I1(1'b0), .CI(n2316), .O(n2314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i15  (.I0(\u_scaler_gray/destx[14] ), 
            .I1(1'b0), .CI(n2321), .O(n2315), .CO(n2316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i14  (.I0(\u_scaler_gray/destx[13] ), 
            .I1(1'b0), .CI(n2323), .O(n2320), .CO(n2321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i13  (.I0(\u_scaler_gray/destx[12] ), 
            .I1(1'b0), .CI(n2325), .O(n2322), .CO(n2323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i12  (.I0(\u_scaler_gray/destx[11] ), 
            .I1(1'b0), .CI(n2327), .O(n2324), .CO(n2325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i11  (.I0(\u_scaler_gray/destx[10] ), 
            .I1(1'b0), .CI(n2329), .O(n2326), .CO(n2327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i10  (.I0(\u_scaler_gray/destx[9] ), 
            .I1(1'b0), .CI(n2331), .O(n2328), .CO(n2329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i9  (.I0(\u_scaler_gray/destx[8] ), 
            .I1(1'b0), .CI(n2335), .O(n2330), .CO(n2331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i8  (.I0(\u_scaler_gray/destx[7] ), 
            .I1(1'b0), .CI(n2337), .O(n2334), .CO(n2335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i7  (.I0(\u_scaler_gray/destx[6] ), 
            .I1(1'b0), .CI(n2339), .O(n2336), .CO(n2337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i6  (.I0(\u_scaler_gray/destx[5] ), 
            .I1(1'b0), .CI(n2344), .O(n2338), .CO(n2339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i5  (.I0(\u_scaler_gray/destx[4] ), 
            .I1(1'b0), .CI(n2347), .O(n2343), .CO(n2344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i4  (.I0(\u_scaler_gray/destx[3] ), 
            .I1(1'b0), .CI(n2353), .O(n2346), .CO(n2347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), .CI(1'b0), 
            .O(n2349), .CO(n2350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_65/i3  (.I0(\u_scaler_gray/destx[2] ), 
            .I1(1'b0), .CI(n917), .O(n2352), .CO(n2353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(192)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_65/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), .CI(n7571), 
            .O(n2355), .CO(n2356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .I1(n5870), .CI(n7572), .CO(n2367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i16  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[15] ), 
            .I1(1'b0), .CI(n2371), .O(n2369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i15  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[14] ), 
            .I1(1'b0), .CI(n2373), .O(n2370), .CO(n2371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i14  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[13] ), 
            .I1(1'b0), .CI(n2375), .O(n2372), .CO(n2373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i13  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[12] ), 
            .I1(1'b0), .CI(n2377), .O(n2374), .CO(n2375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i12  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[11] ), 
            .I1(1'b0), .CI(n2379), .O(n2376), .CO(n2377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i11  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[10] ), 
            .I1(1'b0), .CI(n2381), .O(n2378), .CO(n2379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i10  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[9] ), 
            .I1(1'b0), .CI(n2383), .O(n2380), .CO(n2381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i9  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[8] ), 
            .I1(1'b0), .CI(n2393), .O(n2382), .CO(n2383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i8  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[7] ), 
            .I1(1'b0), .CI(n2395), .O(n2392), .CO(n2393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i7  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[6] ), 
            .I1(1'b0), .CI(n2397), .O(n2394), .CO(n2395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i6  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[5] ), 
            .I1(1'b0), .CI(n2399), .O(n2396), .CO(n2397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i5  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[4] ), 
            .I1(1'b0), .CI(n2401), .O(n2398), .CO(n2399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i4  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[3] ), 
            .I1(1'b0), .CI(n2403), .O(n2400), .CO(n2401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_25/i3  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[2] ), 
            .I1(1'b0), .CI(n912), .O(n2402), .CO(n2403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(91)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_25/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i16  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] ), 
            .I1(1'b0), .CI(n2485), .O(n2483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i15  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] ), 
            .I1(1'b0), .CI(n2487), .O(n2484), .CO(n2485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i14  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] ), 
            .I1(1'b0), .CI(n2489), .O(n2486), .CO(n2487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i13  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] ), 
            .I1(1'b0), .CI(n2491), .O(n2488), .CO(n2489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i12  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] ), 
            .I1(1'b0), .CI(n2493), .O(n2490), .CO(n2491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i11  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] ), 
            .I1(1'b0), .CI(n2495), .O(n2492), .CO(n2493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i10  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] ), 
            .I1(1'b0), .CI(n2497), .O(n2494), .CO(n2495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i9  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] ), 
            .I1(1'b0), .CI(n2499), .O(n2496), .CO(n2497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i8  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] ), 
            .I1(1'b0), .CI(n2523), .O(n2498), .CO(n2499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i3  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(1'b0), .CI(n2513), .O(n2510), .CO(n2511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i2  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), .CI(1'b0), 
            .O(n2512), .CO(n2513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i2  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] ), .CI(1'b0), 
            .O(n2517), .CO(n2518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .CI(n7574), .O(n2520), .CO(n2521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i7  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] ), 
            .I1(1'b0), .CI(n2528), .O(n2522), .CO(n2523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i6  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] ), 
            .I1(1'b0), .CI(n2540), .O(n2527), .CO(n2528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i2  (.I0(\u_lcd_driver/hcnt[1] ), .I1(\u_lcd_driver/hcnt[0] ), 
            .CI(1'b0), .O(n2537), .CO(n2538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(82)
    defparam \u_lcd_driver/add_7/i2 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i5  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] ), 
            .I1(1'b0), .CI(n2542), .O(n2539), .CO(n2540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i4  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] ), 
            .I1(1'b0), .CI(n2544), .O(n2541), .CO(n2542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_16/i3  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] ), 
            .I1(1'b0), .CI(n905), .O(n2543), .CO(n2544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(76)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_16/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i16  (.I0(\u_scaler_gray/vs_cnt[15] ), .I1(1'b0), 
            .CI(n2547), .O(n2545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i15  (.I0(\u_scaler_gray/vs_cnt[14] ), .I1(1'b0), 
            .CI(n2549), .O(n2546), .CO(n2547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i14  (.I0(\u_scaler_gray/vs_cnt[13] ), .I1(1'b0), 
            .CI(n2563), .O(n2548), .CO(n2549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i13  (.I0(\u_scaler_gray/vs_cnt[12] ), .I1(1'b0), 
            .CI(n2565), .O(n2562), .CO(n2563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i12  (.I0(\u_scaler_gray/vs_cnt[11] ), .I1(1'b0), 
            .CI(n2567), .O(n2564), .CO(n2565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i11  (.I0(\u_scaler_gray/vs_cnt[10] ), .I1(1'b0), 
            .CI(n2569), .O(n2566), .CO(n2567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i10  (.I0(\u_scaler_gray/vs_cnt[9] ), .I1(1'b0), 
            .CI(n2571), .O(n2568), .CO(n2569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i9  (.I0(\u_scaler_gray/vs_cnt[8] ), .I1(1'b0), 
            .CI(n2573), .O(n2570), .CO(n2571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i8  (.I0(\u_scaler_gray/vs_cnt[7] ), .I1(1'b0), 
            .CI(n2575), .O(n2572), .CO(n2573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i7  (.I0(\u_scaler_gray/vs_cnt[6] ), .I1(1'b0), 
            .CI(n2577), .O(n2574), .CO(n2575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i6  (.I0(\u_scaler_gray/vs_cnt[5] ), .I1(1'b0), 
            .CI(n2579), .O(n2576), .CO(n2577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i5  (.I0(\u_scaler_gray/vs_cnt[4] ), .I1(1'b0), 
            .CI(n2581), .O(n2578), .CO(n2579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i4  (.I0(\u_scaler_gray/vs_cnt[3] ), .I1(1'b0), 
            .CI(n2583), .O(n2580), .CO(n2581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/add_12/i3  (.I0(\u_scaler_gray/vs_cnt[2] ), .I1(1'b0), 
            .CI(n901), .O(n2582), .CO(n2583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\scaler_gray.v(110)
    defparam \u_scaler_gray/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i16  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15] ), 
            .I1(1'b0), .CI(n2586), .O(n2584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i16 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i15  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14] ), 
            .I1(1'b0), .CI(n2588), .O(n2585), .CO(n2586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i15 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i14  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13] ), 
            .I1(1'b0), .CI(n2590), .O(n2587), .CO(n2588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i14 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i13  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12] ), 
            .I1(1'b0), .CI(n2592), .O(n2589), .CO(n2590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i13 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i12  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11] ), 
            .I1(1'b0), .CI(n2594), .O(n2591), .CO(n2592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i12 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i11  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10] ), 
            .I1(1'b0), .CI(n2596), .O(n2593), .CO(n2594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i11 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i10  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9] ), 
            .I1(1'b0), .CI(n2598), .O(n2595), .CO(n2596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i10 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i9  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8] ), 
            .I1(1'b0), .CI(n2680), .O(n2597), .CO(n2598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i9 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i8  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7] ), 
            .I1(1'b0), .CI(n2682), .O(n2679), .CO(n2680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i8 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i7  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6] ), 
            .I1(1'b0), .CI(n2684), .O(n2681), .CO(n2682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i7 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i6  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5] ), 
            .I1(1'b0), .CI(n2687), .O(n2683), .CO(n2684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i6 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i5  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4] ), 
            .I1(1'b0), .CI(n2691), .O(n2686), .CO(n2687)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i5 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i4  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3] ), 
            .I1(1'b0), .CI(n2693), .O(n2690), .CO(n2691)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i4 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_scaler_gray/u0_data_stream_ctr/add_7/i3  (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2] ), 
            .I1(1'b0), .CI(n736), .O(n2692), .CO(n2693)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\data_stream_ctr.v(60)
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i3 .I0_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/add_7/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i15  (.I0(1'b0), 
            .I1(1'b1), .CI(n2730), .O(n2728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14  (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[13] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] ), 
            .CI(n2732), .O(n2729), .CO(n2730)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13  (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_q ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), .CI(n2734), .O(n2731), 
            .CO(n2732)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12  (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1_q ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[11] ), .CI(n2736), .O(n2733), 
            .CO(n2734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11  (.I0(n6314), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[10] ), .CI(n2738), .O(n2735), 
            .CO(n2736)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10  (.I0(n6317), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[9] ), .CI(n2740), .O(n2737), 
            .CO(n2738)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9  (.I0(n6320), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[8] ), .CI(n2742), .O(n2739), 
            .CO(n2740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8  (.I0(n6323), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[7] ), .CI(n2744), .O(n2741), 
            .CO(n2742)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7  (.I0(n6326), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[6] ), .CI(n2746), .O(n2743), 
            .CO(n2744)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6  (.I0(n6329), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[5] ), .CI(n2748), .O(n2745), 
            .CO(n2746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5  (.I0(n6332), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[4] ), .CI(n2750), .O(n2747), 
            .CO(n2748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4  (.I0(n6335), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[3] ), .CI(n2752), .O(n2749), 
            .CO(n2750)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i3  (.I0(n6338), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[2] ), .CI(n2754), .O(n2751), 
            .CO(n2752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i2  (.I0(n6341), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[1] ), .CI(n722), .O(n2753), 
            .CO(n2754)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1261)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i14  (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] ), 
            .I1(1'b0), .CI(n2757), .O(n2755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i14 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i13  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), 
            .I1(1'b0), .CI(n2759), .O(n2756), .CO(n2757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i13 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i12  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[11] ), 
            .I1(1'b0), .CI(n2761), .O(n2758), .CO(n2759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i12 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i11  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[10] ), 
            .I1(1'b0), .CI(n2763), .O(n2760), .CO(n2761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i11 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i10  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[9] ), 
            .I1(1'b0), .CI(n2765), .O(n2762), .CO(n2763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i10 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[8] ), 
            .I1(1'b0), .CI(n2767), .O(n2764), .CO(n2765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[7] ), 
            .I1(1'b0), .CI(n2769), .O(n2766), .CO(n2767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[6] ), 
            .I1(1'b0), .CI(n2771), .O(n2768), .CO(n2769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[5] ), 
            .I1(1'b0), .CI(n2773), .O(n2770), .CO(n2771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[4] ), 
            .I1(1'b0), .CI(n2775), .O(n2772), .CO(n2773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[3] ), 
            .I1(1'b0), .CI(n2777), .O(n2774), .CO(n2775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3  (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[2] ), 
            .I1(1'b0), .CI(n716), .O(n2776), .CO(n2777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1282)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i14  (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] ), 
            .I1(1'b0), .CI(n2794), .O(n2792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i14 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), 
            .I1(1'b0), .CI(n2796), .O(n2793), .CO(n2794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[11] ), 
            .I1(1'b0), .CI(n2798), .O(n2795), .CO(n2796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[10] ), 
            .I1(1'b0), .CI(n2800), .O(n2797), .CO(n2798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[9] ), 
            .I1(1'b0), .CI(n2802), .O(n2799), .CO(n2800)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[8] ), 
            .I1(1'b0), .CI(n2804), .O(n2801), .CO(n2802)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[7] ), 
            .I1(1'b0), .CI(n2806), .O(n2803), .CO(n2804)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[6] ), 
            .I1(1'b0), .CI(n2808), .O(n2805), .CO(n2806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[5] ), 
            .I1(1'b0), .CI(n2810), .O(n2807), .CO(n2808)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[4] ), 
            .I1(1'b0), .CI(n2812), .O(n2809), .CO(n2810)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4  (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[3] ), 
            .I1(1'b0), .CI(n704), .O(n2811), .CO(n2812)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(1272)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4 .I0_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i9  (.I0(\u_sensor_frame_count/cmos_fps_cnt[8] ), 
            .I1(1'b0), .CI(n2857), .O(n2855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i9 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i8  (.I0(\u_sensor_frame_count/cmos_fps_cnt[7] ), 
            .I1(1'b0), .CI(n2859), .O(n2856), .CO(n2857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i8 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i7  (.I0(\u_sensor_frame_count/cmos_fps_cnt[6] ), 
            .I1(1'b0), .CI(n2861), .O(n2858), .CO(n2859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i7 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i6  (.I0(\u_sensor_frame_count/cmos_fps_cnt[5] ), 
            .I1(1'b0), .CI(n2863), .O(n2860), .CO(n2861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i6 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i5  (.I0(\u_sensor_frame_count/cmos_fps_cnt[4] ), 
            .I1(1'b0), .CI(n2865), .O(n2862), .CO(n2863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i5 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i4  (.I0(\u_sensor_frame_count/cmos_fps_cnt[3] ), 
            .I1(1'b0), .CI(n2867), .O(n2864), .CO(n2865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i4 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_23/i3  (.I0(\u_sensor_frame_count/cmos_fps_cnt[2] ), 
            .I1(1'b0), .CI(n602), .O(n2866), .CO(n2867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(87)
    defparam \u_sensor_frame_count/add_23/i3 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_23/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i28  (.I0(\u_sensor_frame_count/delay_cnt[27] ), 
            .I1(1'b0), .CI(n2870), .O(n2868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i28 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i27  (.I0(\u_sensor_frame_count/delay_cnt[26] ), 
            .I1(1'b0), .CI(n2872), .O(n2869), .CO(n2870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i27 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i26  (.I0(\u_sensor_frame_count/delay_cnt[25] ), 
            .I1(1'b0), .CI(n2874), .O(n2871), .CO(n2872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i26 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i25  (.I0(\u_sensor_frame_count/delay_cnt[24] ), 
            .I1(1'b0), .CI(n2876), .O(n2873), .CO(n2874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i25 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i24  (.I0(\u_sensor_frame_count/delay_cnt[23] ), 
            .I1(1'b0), .CI(n2878), .O(n2875), .CO(n2876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i24 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i23  (.I0(\u_sensor_frame_count/delay_cnt[22] ), 
            .I1(1'b0), .CI(n2880), .O(n2877), .CO(n2878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i23 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i22  (.I0(\u_sensor_frame_count/delay_cnt[21] ), 
            .I1(1'b0), .CI(n2882), .O(n2879), .CO(n2880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i22 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i21  (.I0(\u_sensor_frame_count/delay_cnt[20] ), 
            .I1(1'b0), .CI(n2899), .O(n2881), .CO(n2882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i21 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i20  (.I0(\u_sensor_frame_count/delay_cnt[19] ), 
            .I1(1'b0), .CI(n2901), .O(n2898), .CO(n2899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i20 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i19  (.I0(\u_sensor_frame_count/delay_cnt[18] ), 
            .I1(1'b0), .CI(n3032), .O(n2900), .CO(n2901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i19 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_19/i2  (.I0(\u_lcd_driver/vcnt[1] ), .I1(\u_lcd_driver/vcnt[0] ), 
            .CI(1'b0), .O(n3029), .CO(n3030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(102)
    defparam \u_lcd_driver/add_19/i2 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_19/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i18  (.I0(\u_sensor_frame_count/delay_cnt[17] ), 
            .I1(1'b0), .CI(n3036), .O(n3031), .CO(n3032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i18 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i17  (.I0(\u_sensor_frame_count/delay_cnt[16] ), 
            .I1(1'b0), .CI(n3038), .O(n3035), .CO(n3036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i17 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i16  (.I0(\u_sensor_frame_count/delay_cnt[15] ), 
            .I1(1'b0), .CI(n3042), .O(n3037), .CO(n3038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i16 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_75/i2  (.I0(n362), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .CI(1'b0), .O(n3039), .CO(n3040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(88)
    defparam \u_rgb2dvi/enc_0/add_75/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_75/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_sensor_frame_count/add_14/i15  (.I0(\u_sensor_frame_count/delay_cnt[14] ), 
            .I1(1'b0), .CI(n3046), .O(n3041), .CO(n3042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i15 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i14  (.I0(\u_sensor_frame_count/delay_cnt[13] ), 
            .I1(1'b0), .CI(n3048), .O(n3045), .CO(n3046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i14 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i13  (.I0(\u_sensor_frame_count/delay_cnt[12] ), 
            .I1(1'b0), .CI(n3053), .O(n3047), .CO(n3048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i13 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i12  (.I0(\u_sensor_frame_count/delay_cnt[11] ), 
            .I1(1'b0), .CI(n3055), .O(n3052), .CO(n3053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i12 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i11  (.I0(\u_sensor_frame_count/delay_cnt[10] ), 
            .I1(1'b0), .CI(n3068), .O(n3054), .CO(n3055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i11 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i10  (.I0(\u_sensor_frame_count/delay_cnt[9] ), 
            .I1(1'b0), .CI(n3070), .O(n3067), .CO(n3068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i10 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i9  (.I0(\u_sensor_frame_count/delay_cnt[8] ), 
            .I1(1'b0), .CI(n3072), .O(n3069), .CO(n3070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i9 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i8  (.I0(\u_sensor_frame_count/delay_cnt[7] ), 
            .I1(1'b0), .CI(n3074), .O(n3071), .CO(n3072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i8 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i7  (.I0(\u_sensor_frame_count/delay_cnt[6] ), 
            .I1(1'b0), .CI(n3076), .O(n3073), .CO(n3074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i7 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i6  (.I0(\u_sensor_frame_count/delay_cnt[5] ), 
            .I1(1'b0), .CI(n3078), .O(n3075), .CO(n3076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i6 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i5  (.I0(\u_sensor_frame_count/delay_cnt[4] ), 
            .I1(1'b0), .CI(n3080), .O(n3077), .CO(n3078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i5 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i4  (.I0(\u_sensor_frame_count/delay_cnt[3] ), 
            .I1(1'b0), .CI(n3082), .O(n3079), .CO(n3080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i4 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_sensor_frame_count/add_14/i3  (.I0(\u_sensor_frame_count/delay_cnt[2] ), 
            .I1(1'b0), .CI(n576), .O(n3081), .CO(n3082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\sensor_frame_count.v(69)
    defparam \u_sensor_frame_count/add_14/i3 .I0_POLARITY = 1'b1;
    defparam \u_sensor_frame_count/add_14/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/add_105/i1  (.I0(\u_rgb2dvi/enc_0/acc[0] ), .I1(n3335), 
            .CI(1'b0), .O(n3195), .CO(n3196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_0/add_105/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/add_105/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_0/sub_79/add_2/i2  (.I0(n369), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .CI(n7575), .O(n3207), .CO(n3208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(93)
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_0/sub_79/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i12  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[11] ), 
            .I1(1'b0), .CI(n3211), .O(n3209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i12 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i11  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[10] ), 
            .I1(1'b0), .CI(n3213), .O(n3210), .CO(n3211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i11 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i10  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[9] ), 
            .I1(1'b0), .CI(n3215), .O(n3212), .CO(n3213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i10 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i9  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[8] ), 
            .I1(1'b0), .CI(n3217), .O(n3214), .CO(n3215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i9 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i8  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[7] ), 
            .I1(1'b0), .CI(n3219), .O(n3216), .CO(n3217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i8 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i7  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[6] ), 
            .I1(1'b0), .CI(n3221), .O(n3218), .CO(n3219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i7 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i6  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[5] ), 
            .I1(1'b0), .CI(n3223), .O(n3220), .CO(n3221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i6 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i5  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[4] ), 
            .I1(1'b0), .CI(n3225), .O(n3222), .CO(n3223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i5 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i4  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[3] ), 
            .I1(1'b0), .CI(n3227), .O(n3224), .CO(n3225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i4 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_CMOS_Capture_RAW_Gray/add_30/i3  (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[2] ), 
            .I1(1'b0), .CI(n444), .O(n3226), .CO(n3227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\CMOS_Capture_RAW_Gray.v(106)
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i3 .I0_POLARITY = 1'b1;
    defparam \u_CMOS_Capture_RAW_Gray/add_30/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_1/add_105/i1  (.I0(\u_rgb2dvi/enc_1/acc[0] ), .I1(n3335), 
            .CI(1'b0), .O(n3254), .CO(n3255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_1/add_105/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_1/add_105/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i8  (.I0(\i2c_config_index[7] ), 
            .I1(1'b0), .CI(n3286), .O(n3284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i8 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i7  (.I0(\i2c_config_index[6] ), 
            .I1(1'b0), .CI(n3288), .O(n3285), .CO(n3286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i7 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i6  (.I0(\i2c_config_index[5] ), 
            .I1(1'b0), .CI(n3290), .O(n3287), .CO(n3288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i6 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i5  (.I0(\i2c_config_index[4] ), 
            .I1(1'b0), .CI(n3292), .O(n3289), .CO(n3290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i5 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i4  (.I0(\i2c_config_index[3] ), 
            .I1(1'b0), .CI(n3294), .O(n3291), .CO(n3292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i4 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_50/i3  (.I0(\i2c_config_index[2] ), 
            .I1(1'b0), .CI(n223), .O(n3293), .CO(n3294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(188)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i3 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_50/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i16  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15] ), 
            .I1(1'b0), .CI(n3297), .O(n3295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i16 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i15  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14] ), 
            .I1(1'b0), .CI(n3299), .O(n3296), .CO(n3297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i15 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i14  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13] ), 
            .I1(1'b0), .CI(n3310), .O(n3298), .CO(n3299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i14 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i13  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), 
            .I1(1'b0), .CI(n3312), .O(n3309), .CO(n3310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i13 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i12  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] ), 
            .I1(1'b0), .CI(n3314), .O(n3311), .CO(n3312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i12 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i11  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), 
            .I1(1'b0), .CI(n3316), .O(n3313), .CO(n3314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i11 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i10  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), 
            .I1(1'b0), .CI(n3322), .O(n3315), .CO(n3316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i10 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i9  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] ), 
            .I1(1'b0), .CI(n3324), .O(n3321), .CO(n3322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i9 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i8  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), 
            .I1(1'b0), .CI(n3326), .O(n3323), .CO(n3324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i8 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i7  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] ), 
            .I1(1'b0), .CI(n3328), .O(n3325), .CO(n3326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i7 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i6  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] ), 
            .I1(1'b0), .CI(n3330), .O(n3327), .CO(n3328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i6 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i5  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4] ), 
            .I1(1'b0), .CI(n3334), .O(n3329), .CO(n3330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i5 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/add_105/i1  (.I0(\u_rgb2dvi/enc_2/acc[0] ), .I1(n3335), 
            .CI(1'b0), .O(n3331), .CO(n3332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(98)
    defparam \u_rgb2dvi/enc_2/add_105/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/add_105/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i4  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3] ), 
            .I1(1'b0), .CI(n3339), .O(n3333), .CO(n3334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i4 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_rgb2dvi/enc_2/sub_50/add_2/i1  (.I0(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q ), .CI(n7576), 
            .O(n3335), .CO(n7577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\hdmi_ip\tmds_channel.v(74)
    defparam \u_rgb2dvi/enc_2/sub_50/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_rgb2dvi/enc_2/sub_50/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_16/i3  (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2] ), 
            .I1(1'b0), .CI(n220), .O(n3338), .CO(n3339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(104)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i3 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_16/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i20  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19] ), 
            .I1(1'b0), .CI(n3343), .O(n3341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i20 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i19  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18] ), 
            .I1(1'b0), .CI(n3345), .O(n3342), .CO(n3343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i19 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i18  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17] ), 
            .I1(1'b0), .CI(n3347), .O(n3344), .CO(n3345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i18 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i17  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16] ), 
            .I1(1'b0), .CI(n3349), .O(n3346), .CO(n3347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i17 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i16  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15] ), 
            .I1(1'b0), .CI(n3351), .O(n3348), .CO(n3349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i16 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i15  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14] ), 
            .I1(1'b0), .CI(n3353), .O(n3350), .CO(n3351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i15 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i14  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13] ), 
            .I1(1'b0), .CI(n3355), .O(n3352), .CO(n3353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i14 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i13  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12] ), 
            .I1(1'b0), .CI(n3357), .O(n3354), .CO(n3355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i13 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i12  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11] ), 
            .I1(1'b0), .CI(n3359), .O(n3356), .CO(n3357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i12 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i11  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10] ), 
            .I1(1'b0), .CI(n3361), .O(n3358), .CO(n3359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i11 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i10  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9] ), 
            .I1(1'b0), .CI(n3371), .O(n3360), .CO(n3361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i10 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i9  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8] ), 
            .I1(1'b0), .CI(n3373), .O(n3370), .CO(n3371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i9 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i8  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7] ), 
            .I1(1'b0), .CI(n3375), .O(n3372), .CO(n3373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i8 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i7  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6] ), 
            .I1(1'b0), .CI(n3377), .O(n3374), .CO(n3375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i7 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i6  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5] ), 
            .I1(1'b0), .CI(n3379), .O(n3376), .CO(n3377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i6 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i5  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4] ), 
            .I1(1'b0), .CI(n3381), .O(n3378), .CO(n3379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i5 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i4  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3] ), 
            .I1(1'b0), .CI(n3383), .O(n3380), .CO(n3381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i4 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_i2c_timing_ctrl_16reg_16bit/add_7/i3  (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2] ), 
            .I1(1'b0), .CI(n198), .O(n3382), .CO(n3383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\cmos_i2c\i2c_timing_ctrl_reg16_dat16.v(69)
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i3 .I0_POLARITY = 1'b1;
    defparam \u_i2c_timing_ctrl_16reg_16bit/add_7/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] ), 
            .I1(1'b1), .CI(n3390), .O(n3388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] ), 
            .I1(1'b1), .CI(n3392), .O(n3389), .CO(n3390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] ), 
            .I1(1'b1), .CI(n3394), .O(n3391), .CO(n3392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] ), 
            .I1(1'b1), .CI(n3396), .O(n3393), .CO(n3394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] ), 
            .I1(1'b1), .CI(n3398), .O(n3395), .CO(n3396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] ), 
            .I1(1'b1), .CI(n3400), .O(n3397), .CO(n3398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] ), 
            .I1(1'b1), .CI(n3402), .O(n3399), .CO(n3400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] ), 
            .I1(1'b1), .CI(n3404), .O(n3401), .CO(n3402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] ), 
            .I1(1'b1), .CI(n3406), .O(n3403), .CO(n3404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] ), 
            .I1(1'b1), .CI(n3408), .O(n3405), .CO(n3406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] ), 
            .I1(1'b1), .CI(n3410), .O(n3407), .CO(n3408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] ), 
            .I1(1'b1), .CI(n3412), .O(n3409), .CO(n3410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] ), 
            .I1(1'b1), .CI(n3414), .O(n3411), .CO(n3412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] ), 
            .I1(1'b1), .CI(n3416), .O(n3413), .CO(n3414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] ), 
            .I1(1'b1), .CI(n3418), .O(n3415), .CO(n3416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] ), 
            .I1(1'b1), .CI(n3420), .O(n3417), .CO(n3418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] ), 
            .I1(1'b1), .CI(n3422), .O(n3419), .CO(n3420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] ), 
            .I1(1'b1), .CI(n3424), .O(n3421), .CO(n3422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] ), 
            .I1(1'b1), .CI(n177), .O(n3423), .CO(n3424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i8  (.I0(\PowerOnResetCnt[7] ), .I1(1'b0), .CI(n3428), 
            .O(n3426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i8 .I0_POLARITY = 1'b1;
    defparam \add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i7  (.I0(\PowerOnResetCnt[6] ), .I1(1'b0), .CI(n3430), 
            .O(n3427), .CO(n3428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i7 .I0_POLARITY = 1'b1;
    defparam \add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i6  (.I0(\PowerOnResetCnt[5] ), .I1(1'b0), .CI(n3466), 
            .O(n3429), .CO(n3430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i6 .I0_POLARITY = 1'b1;
    defparam \add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i5  (.I0(\PowerOnResetCnt[4] ), .I1(1'b0), .CI(n3468), 
            .O(n3465), .CO(n3466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i5 .I0_POLARITY = 1'b1;
    defparam \add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i4  (.I0(\PowerOnResetCnt[3] ), .I1(1'b0), .CI(n3470), 
            .O(n3467), .CO(n3468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i4 .I0_POLARITY = 1'b1;
    defparam \add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i3  (.I0(\PowerOnResetCnt[2] ), .I1(1'b0), .CI(n3472), 
            .O(n3469), .CO(n3470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i3 .I0_POLARITY = 1'b1;
    defparam \add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i2  (.I0(\PowerOnResetCnt[1] ), .I1(1'b0), .CI(n3474), 
            .O(n3471), .CO(n3472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i2 .I0_POLARITY = 1'b1;
    defparam \add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_10/i1  (.I0(\PowerOnResetCnt[0] ), .I1(\reduce_nand_9/n7 ), 
            .CI(1'b0), .O(n3473), .CO(n3474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\T35_Sensor_DDR3_LCD_Test.v(120)
    defparam \add_10/i1 .I0_POLARITY = 1'b1;
    defparam \add_10/i1 .I1_POLARITY = 1'b0;
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2105_2), .WDATA({\cmos_frame_Gray[2] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n98 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3b12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2091_2), .WDATA({\cmos_frame_Gray[0] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n105 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$02 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2091_2), .WDATA({\cmos_frame_Gray[2] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n99 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0b12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2091_2), .WDATA({\cmos_frame_Gray[1] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n102 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$012 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2105_2), .WDATA({\cmos_frame_Gray[0] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n104 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$32 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2091_2), .WDATA({\cmos_frame_Gray[3] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n96 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0c12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2091_2), .WDATA({\cmos_frame_Gray[4] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n93 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0d12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2091_2), .WDATA({\cmos_frame_Gray[5] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n90 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0e12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2091_2), .WDATA({\cmos_frame_Gray[6] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n87 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0f12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 ), 
            .RE(n2091_2), .WDATA({\cmos_frame_Gray[7] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n84 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$0g1 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2105_2), .WDATA({\cmos_frame_Gray[1] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n101 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$312 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2105_2), .WDATA({\cmos_frame_Gray[3] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n95 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3c12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2105_2), .WDATA({\cmos_frame_Gray[4] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n92 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3d12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2105_2), .WDATA({\cmos_frame_Gray[5] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n89 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3e12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2105_2), .WDATA({\cmos_frame_Gray[6] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n86 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3f12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1  (.WCLK(\cmos_pclk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 ), 
            .RE(n2105_2), .WDATA({\cmos_frame_Gray[7] }), .WADDR({\u_afifo_buf/u_efx_fifo_top/waddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[10] , \u_afifo_buf/u_efx_fifo_top/waddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[8] , \u_afifo_buf/u_efx_fifo_top/waddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[6] , \u_afifo_buf/u_efx_fifo_top/waddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[4] , \u_afifo_buf/u_efx_fifo_top/waddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[2] , \u_afifo_buf/u_efx_fifo_top/waddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/waddr[0] }), .RADDR({\u_afifo_buf/u_efx_fifo_top/raddr[11] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[10] , \u_afifo_buf/u_efx_fifo_top/raddr[9] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[8] , \u_afifo_buf/u_efx_fifo_top/raddr[7] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[6] , \u_afifo_buf/u_efx_fifo_top/raddr[5] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[4] , \u_afifo_buf/u_efx_fifo_top/raddr[3] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[2] , \u_afifo_buf/u_efx_fifo_top/raddr[1] , 
            \u_afifo_buf/u_efx_fifo_top/raddr[0] }), .RDATA({\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n83 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(705)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .READ_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .WRITE_WIDTH = 1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .WCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .WE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .RCLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .RE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .OUTPUT_REG = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/ram__D$3g1 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[6] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_1=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_2=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_3=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_4=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_5=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_6=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_7=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_0 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_1 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_2 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_3 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_4 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_5 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_6 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_7 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[1] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_1=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_2=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_3=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_4=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_5=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_6=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_7=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_0 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_1 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_2 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_3 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_4 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_5 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_6 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_7 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[1] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_1=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_2=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_3=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_4=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_5=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_6=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_7=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_0 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_1 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_2 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_3 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_4 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_5 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_6 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_7 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[1] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_1=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_2=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_3=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_4=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_5=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_6=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_7=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_0 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_1 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_2 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_3 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_4 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_5 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_6 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_7 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[1] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_1=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_2=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_3=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_4=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_5=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_6=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_7=256'h3333333333333333333333333333333333333333333333333333333333333333, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_0 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_1 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_2 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_3 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_4 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_5 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_6 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_7 = 256'h3333333333333333333333333333333333333333333333333333333333333333;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[5] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_1=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_2=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_3=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_4=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_5=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_6=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_7=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_0 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_1 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_2 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_3 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_4 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_5 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_6 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_7 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[7] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_1=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_2=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_3=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_4=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_5=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_6=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_7=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_0 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_1 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_2 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_3 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_4 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_5 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_6 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_7 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[4] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_1=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_2=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_3=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_4=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_5=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_6=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_7=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_0 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_1 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_2 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_3 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_4 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_5 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_6 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_7 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[2] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_1=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_2=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_3=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_4=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_5=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_6=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_7=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_0 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_1 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_2 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_3 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_4 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_5 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_6 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_7 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[3] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_1=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_2=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_3=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_4=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_5=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_6=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_7=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_0 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_1 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_2 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_3 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_4 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_5 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_6 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_7 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[6] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_1=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_2=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_3=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_4=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_5=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_6=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_7=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_0 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_1 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_2 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_3 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_4 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_5 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_6 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_7 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[0] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata00[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_1=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_2=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_3=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_4=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_5=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_6=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_7=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_0 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_1 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_2 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_3 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_4 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_5 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_6 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_7 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram00/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[5] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_1=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_2=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_3=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_4=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_5=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_6=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_7=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_0 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_1 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_2 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_3 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_4 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_5 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_6 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_7 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[7] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_1=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_2=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_3=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_4=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_5=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_6=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_7=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_0 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_1 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_2 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_3 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_4 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_5 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_6 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_7 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[4] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_1=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_2=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_3=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_4=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_5=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_6=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_7=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_0 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_1 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_2 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_3 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_4 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_5 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_6 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_7 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[2] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_1=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_2=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_3=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_4=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_5=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_6=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_7=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_0 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_1 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_2 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_3 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_4 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_5 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_6 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_7 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[3] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_1=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_2=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_3=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_4=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_5=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_6=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_7=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_0 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_1 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_2 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_3 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_4 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_5 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_6 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_7 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[6] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_1=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_2=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_3=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_4=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_5=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_6=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_7=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_0 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_1 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_2 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_3 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_4 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_5 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_6 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_7 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[0] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata01[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_1=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_2=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_3=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_4=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_5=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_6=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_7=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_0 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_1 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_2 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_3 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_4 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_5 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_6 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_7 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram01/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[5] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_1=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_2=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_3=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_4=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_5=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_6=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_7=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_0 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_1 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_2 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_3 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_4 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_5 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_6 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_7 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[7] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_1=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_2=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_3=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_4=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_5=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_6=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_7=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_0 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_1 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_2 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_3 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_4 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_5 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_6 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_7 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[4] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_1=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_2=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_3=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_4=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_5=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_6=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_7=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_0 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_1 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_2 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_3 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_4 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_5 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_6 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_7 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[2] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_1=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_2=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_3=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_4=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_5=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_6=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_7=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_0 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_1 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_2 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_3 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_4 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_5 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_6 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_7 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[3] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_1=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_2=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_3=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_4=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_5=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_6=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_7=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_0 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_1 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_2 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_3 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_4 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_5 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_6 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_7 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[6] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_1=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_2=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_3=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_4=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_5=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_6=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_7=256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_0 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_1 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_2 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_3 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_4 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_5 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_6 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_7 = 256'h0000000000000000FFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[0] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I }), .RDATA({\u_scaler_gray/tdata10[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_1=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_2=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_3=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_4=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_5=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_6=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_7=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_0 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_1 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_2 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_3 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_4 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_5 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_6 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_7 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram10/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[5] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_1=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_2=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_3=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_4=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_5=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_6=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_7=256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_0 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_1 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_2 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_3 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_4 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_5 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_6 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_7 = 256'h00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF00000000FFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[7] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_1=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_2=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_3=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_4=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_5=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_6=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_7=256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_0 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_1 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_2 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_3 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_4 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_5 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_6 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_7 = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[4] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_1=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_2=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_3=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_4=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_5=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_6=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_7=256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_0 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_1 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_2 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_3 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_4 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_5 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_6 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_7 = 256'h0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF0000FFFF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[2] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_1=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_2=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_3=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_4=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_5=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_6=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_7=256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_0 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_1 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_2 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_3 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_4 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_5 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_6 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_7 = 256'h0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[3] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_1=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_2=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_3=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_4=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_5=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_6=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_7=256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_0 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_1 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_2 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_3 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_4 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_5 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_6 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_7 = 256'h00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF00FF;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(n197_2), .RE(\u_scaler_gray/u0_data_stream_ctr/scaler_valid_d[3] ), 
            .WDATA({\tdata_i[0] }), .WADDR({\u_scaler_gray/u0_data_stream_ctr/w_addra[11] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[10] , \u_scaler_gray/u0_data_stream_ctr/w_addra[9] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[8] , \u_scaler_gray/u0_data_stream_ctr/w_addra[7] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[6] , \u_scaler_gray/u0_data_stream_ctr/w_addra[5] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[4] , \u_scaler_gray/u0_data_stream_ctr/w_addra[3] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[2] , \u_scaler_gray/u0_data_stream_ctr/w_addra[1] , 
            \u_scaler_gray/u0_data_stream_ctr/w_addra[0] }), .RADDR({\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I , \u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I , 
            \u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I }), .RDATA({\u_scaler_gray/tdata11[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_1=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_2=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_3=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_4=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_5=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_6=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_7=256'h5555555555555555555555555555555555555555555555555555555555555555, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\simple_dual_port_ram.v(19)
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .READ_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_0 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_1 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_2 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_3 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_4 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_5 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_6 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_7 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .OUTPUT_REG = 1'b1;
    defparam \u_scaler_gray/u0_data_stream_ctr/u_simple_dual_port_ram11/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[4] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[4], DdrCtrl_WDATA_0[12], DdrCtrl_WDATA_0[20], 
            DdrCtrl_WDATA_0[28], DdrCtrl_WDATA_0[36], DdrCtrl_WDATA_0[44], 
            DdrCtrl_WDATA_0[52], DdrCtrl_WDATA_0[60], DdrCtrl_WDATA_0[68], 
            DdrCtrl_WDATA_0[76], DdrCtrl_WDATA_0[84], DdrCtrl_WDATA_0[92], 
            DdrCtrl_WDATA_0[100], DdrCtrl_WDATA_0[108], DdrCtrl_WDATA_0[116], 
            DdrCtrl_WDATA_0[124]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[1] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[1], DdrCtrl_WDATA_0[9], DdrCtrl_WDATA_0[17], 
            DdrCtrl_WDATA_0[25], DdrCtrl_WDATA_0[33], DdrCtrl_WDATA_0[41], 
            DdrCtrl_WDATA_0[49], DdrCtrl_WDATA_0[57], DdrCtrl_WDATA_0[65], 
            DdrCtrl_WDATA_0[73], DdrCtrl_WDATA_0[81], DdrCtrl_WDATA_0[89], 
            DdrCtrl_WDATA_0[97], DdrCtrl_WDATA_0[105], DdrCtrl_WDATA_0[113], 
            DdrCtrl_WDATA_0[121]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[0] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[0], DdrCtrl_WDATA_0[8], DdrCtrl_WDATA_0[16], 
            DdrCtrl_WDATA_0[24], DdrCtrl_WDATA_0[32], DdrCtrl_WDATA_0[40], 
            DdrCtrl_WDATA_0[48], DdrCtrl_WDATA_0[56], DdrCtrl_WDATA_0[64], 
            DdrCtrl_WDATA_0[72], DdrCtrl_WDATA_0[80], DdrCtrl_WDATA_0[88], 
            DdrCtrl_WDATA_0[96], DdrCtrl_WDATA_0[104], DdrCtrl_WDATA_0[112], 
            DdrCtrl_WDATA_0[120]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[2] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[2], DdrCtrl_WDATA_0[10], DdrCtrl_WDATA_0[18], 
            DdrCtrl_WDATA_0[26], DdrCtrl_WDATA_0[34], DdrCtrl_WDATA_0[42], 
            DdrCtrl_WDATA_0[50], DdrCtrl_WDATA_0[58], DdrCtrl_WDATA_0[66], 
            DdrCtrl_WDATA_0[74], DdrCtrl_WDATA_0[82], DdrCtrl_WDATA_0[90], 
            DdrCtrl_WDATA_0[98], DdrCtrl_WDATA_0[106], DdrCtrl_WDATA_0[114], 
            DdrCtrl_WDATA_0[122]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[5] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[5], DdrCtrl_WDATA_0[13], DdrCtrl_WDATA_0[21], 
            DdrCtrl_WDATA_0[29], DdrCtrl_WDATA_0[37], DdrCtrl_WDATA_0[45], 
            DdrCtrl_WDATA_0[53], DdrCtrl_WDATA_0[61], DdrCtrl_WDATA_0[69], 
            DdrCtrl_WDATA_0[77], DdrCtrl_WDATA_0[85], DdrCtrl_WDATA_0[93], 
            DdrCtrl_WDATA_0[101], DdrCtrl_WDATA_0[109], DdrCtrl_WDATA_0[117], 
            DdrCtrl_WDATA_0[125]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[7] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[7], DdrCtrl_WDATA_0[15], DdrCtrl_WDATA_0[23], 
            DdrCtrl_WDATA_0[31], DdrCtrl_WDATA_0[39], DdrCtrl_WDATA_0[47], 
            DdrCtrl_WDATA_0[55], DdrCtrl_WDATA_0[63], DdrCtrl_WDATA_0[71], 
            DdrCtrl_WDATA_0[79], DdrCtrl_WDATA_0[87], DdrCtrl_WDATA_0[95], 
            DdrCtrl_WDATA_0[103], DdrCtrl_WDATA_0[111], DdrCtrl_WDATA_0[119], 
            DdrCtrl_WDATA_0[127]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[6] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[6], DdrCtrl_WDATA_0[14], DdrCtrl_WDATA_0[22], 
            DdrCtrl_WDATA_0[30], DdrCtrl_WDATA_0[38], DdrCtrl_WDATA_0[46], 
            DdrCtrl_WDATA_0[54], DdrCtrl_WDATA_0[62], DdrCtrl_WDATA_0[70], 
            DdrCtrl_WDATA_0[78], DdrCtrl_WDATA_0[86], DdrCtrl_WDATA_0[94], 
            DdrCtrl_WDATA_0[102], DdrCtrl_WDATA_0[110], DdrCtrl_WDATA_0[118], 
            DdrCtrl_WDATA_0[126]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[1] , 
            \u_axi4_ctrl/rfifo_wdata[9] , \u_axi4_ctrl/rfifo_wdata[17] , 
            \u_axi4_ctrl/rfifo_wdata[25] , \u_axi4_ctrl/rfifo_wdata[33] , 
            \u_axi4_ctrl/rfifo_wdata[41] , \u_axi4_ctrl/rfifo_wdata[49] , 
            \u_axi4_ctrl/rfifo_wdata[57] , \u_axi4_ctrl/rfifo_wdata[65] , 
            \u_axi4_ctrl/rfifo_wdata[73] , \u_axi4_ctrl/rfifo_wdata[81] , 
            \u_axi4_ctrl/rfifo_wdata[89] , \u_axi4_ctrl/rfifo_wdata[97] , 
            \u_axi4_ctrl/rfifo_wdata[105] , \u_axi4_ctrl/rfifo_wdata[113] , 
            \u_axi4_ctrl/rfifo_wdata[121] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[1] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\tdata_o[3] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({DdrCtrl_WDATA_0[3], DdrCtrl_WDATA_0[11], DdrCtrl_WDATA_0[19], 
            DdrCtrl_WDATA_0[27], DdrCtrl_WDATA_0[35], DdrCtrl_WDATA_0[43], 
            DdrCtrl_WDATA_0[51], DdrCtrl_WDATA_0[59], DdrCtrl_WDATA_0[67], 
            DdrCtrl_WDATA_0[75], DdrCtrl_WDATA_0[83], DdrCtrl_WDATA_0[91], 
            DdrCtrl_WDATA_0[99], DdrCtrl_WDATA_0[107], DdrCtrl_WDATA_0[115], 
            DdrCtrl_WDATA_0[123]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=16, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .READ_WIDTH = 16;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[5] , 
            \u_axi4_ctrl/rfifo_wdata[13] , \u_axi4_ctrl/rfifo_wdata[21] , 
            \u_axi4_ctrl/rfifo_wdata[29] , \u_axi4_ctrl/rfifo_wdata[37] , 
            \u_axi4_ctrl/rfifo_wdata[45] , \u_axi4_ctrl/rfifo_wdata[53] , 
            \u_axi4_ctrl/rfifo_wdata[61] , \u_axi4_ctrl/rfifo_wdata[69] , 
            \u_axi4_ctrl/rfifo_wdata[77] , \u_axi4_ctrl/rfifo_wdata[85] , 
            \u_axi4_ctrl/rfifo_wdata[93] , \u_axi4_ctrl/rfifo_wdata[101] , 
            \u_axi4_ctrl/rfifo_wdata[109] , \u_axi4_ctrl/rfifo_wdata[117] , 
            \u_axi4_ctrl/rfifo_wdata[125] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[5] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[3] , 
            \u_axi4_ctrl/rfifo_wdata[11] , \u_axi4_ctrl/rfifo_wdata[19] , 
            \u_axi4_ctrl/rfifo_wdata[27] , \u_axi4_ctrl/rfifo_wdata[35] , 
            \u_axi4_ctrl/rfifo_wdata[43] , \u_axi4_ctrl/rfifo_wdata[51] , 
            \u_axi4_ctrl/rfifo_wdata[59] , \u_axi4_ctrl/rfifo_wdata[67] , 
            \u_axi4_ctrl/rfifo_wdata[75] , \u_axi4_ctrl/rfifo_wdata[83] , 
            \u_axi4_ctrl/rfifo_wdata[91] , \u_axi4_ctrl/rfifo_wdata[99] , 
            \u_axi4_ctrl/rfifo_wdata[107] , \u_axi4_ctrl/rfifo_wdata[115] , 
            \u_axi4_ctrl/rfifo_wdata[123] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[3] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[7] , 
            \u_axi4_ctrl/rfifo_wdata[15] , \u_axi4_ctrl/rfifo_wdata[23] , 
            \u_axi4_ctrl/rfifo_wdata[31] , \u_axi4_ctrl/rfifo_wdata[39] , 
            \u_axi4_ctrl/rfifo_wdata[47] , \u_axi4_ctrl/rfifo_wdata[55] , 
            \u_axi4_ctrl/rfifo_wdata[63] , \u_axi4_ctrl/rfifo_wdata[71] , 
            \u_axi4_ctrl/rfifo_wdata[79] , \u_axi4_ctrl/rfifo_wdata[87] , 
            \u_axi4_ctrl/rfifo_wdata[95] , \u_axi4_ctrl/rfifo_wdata[103] , 
            \u_axi4_ctrl/rfifo_wdata[111] , \u_axi4_ctrl/rfifo_wdata[119] , 
            \u_axi4_ctrl/rfifo_wdata[127] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[7] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[2] , 
            \u_axi4_ctrl/rfifo_wdata[10] , \u_axi4_ctrl/rfifo_wdata[18] , 
            \u_axi4_ctrl/rfifo_wdata[26] , \u_axi4_ctrl/rfifo_wdata[34] , 
            \u_axi4_ctrl/rfifo_wdata[42] , \u_axi4_ctrl/rfifo_wdata[50] , 
            \u_axi4_ctrl/rfifo_wdata[58] , \u_axi4_ctrl/rfifo_wdata[66] , 
            \u_axi4_ctrl/rfifo_wdata[74] , \u_axi4_ctrl/rfifo_wdata[82] , 
            \u_axi4_ctrl/rfifo_wdata[90] , \u_axi4_ctrl/rfifo_wdata[98] , 
            \u_axi4_ctrl/rfifo_wdata[106] , \u_axi4_ctrl/rfifo_wdata[114] , 
            \u_axi4_ctrl/rfifo_wdata[122] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[6] , 
            \u_axi4_ctrl/rfifo_wdata[14] , \u_axi4_ctrl/rfifo_wdata[22] , 
            \u_axi4_ctrl/rfifo_wdata[30] , \u_axi4_ctrl/rfifo_wdata[38] , 
            \u_axi4_ctrl/rfifo_wdata[46] , \u_axi4_ctrl/rfifo_wdata[54] , 
            \u_axi4_ctrl/rfifo_wdata[62] , \u_axi4_ctrl/rfifo_wdata[70] , 
            \u_axi4_ctrl/rfifo_wdata[78] , \u_axi4_ctrl/rfifo_wdata[86] , 
            \u_axi4_ctrl/rfifo_wdata[94] , \u_axi4_ctrl/rfifo_wdata[102] , 
            \u_axi4_ctrl/rfifo_wdata[110] , \u_axi4_ctrl/rfifo_wdata[118] , 
            \u_axi4_ctrl/rfifo_wdata[126] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[0] , 
            \u_axi4_ctrl/rfifo_wdata[8] , \u_axi4_ctrl/rfifo_wdata[16] , 
            \u_axi4_ctrl/rfifo_wdata[24] , \u_axi4_ctrl/rfifo_wdata[32] , 
            \u_axi4_ctrl/rfifo_wdata[40] , \u_axi4_ctrl/rfifo_wdata[48] , 
            \u_axi4_ctrl/rfifo_wdata[56] , \u_axi4_ctrl/rfifo_wdata[64] , 
            \u_axi4_ctrl/rfifo_wdata[72] , \u_axi4_ctrl/rfifo_wdata[80] , 
            \u_axi4_ctrl/rfifo_wdata[88] , \u_axi4_ctrl/rfifo_wdata[96] , 
            \u_axi4_ctrl/rfifo_wdata[104] , \u_axi4_ctrl/rfifo_wdata[112] , 
            \u_axi4_ctrl/rfifo_wdata[120] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\hdmi_clk1x_i~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[4] , 
            \u_axi4_ctrl/rfifo_wdata[12] , \u_axi4_ctrl/rfifo_wdata[20] , 
            \u_axi4_ctrl/rfifo_wdata[28] , \u_axi4_ctrl/rfifo_wdata[36] , 
            \u_axi4_ctrl/rfifo_wdata[44] , \u_axi4_ctrl/rfifo_wdata[52] , 
            \u_axi4_ctrl/rfifo_wdata[60] , \u_axi4_ctrl/rfifo_wdata[68] , 
            \u_axi4_ctrl/rfifo_wdata[76] , \u_axi4_ctrl/rfifo_wdata[84] , 
            \u_axi4_ctrl/rfifo_wdata[92] , \u_axi4_ctrl/rfifo_wdata[100] , 
            \u_axi4_ctrl/rfifo_wdata[108] , \u_axi4_ctrl/rfifo_wdata[116] , 
            \u_axi4_ctrl/rfifo_wdata[124] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({\lcd_data[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .READ_WIDTH = 1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, n1163, n1164, n1166, n1168, 
            n1170, n1172, n1174, n1176, n1178, n1180, n1182, n1719}), 
            .B({10'b0000000000, \u_scaler_gray/tdata01[7] , \u_scaler_gray/tdata01[6] , 
            \u_scaler_gray/tdata01[5] , \u_scaler_gray/tdata01[4] , \u_scaler_gray/tdata01[3] , 
            \u_scaler_gray/tdata01[2] , \u_scaler_gray/tdata01[1] , \u_scaler_gray/tdata01[0] }), 
            .O({Open_0, Open_1, Open_2, Open_3, Open_4, Open_5, 
            Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, Open_12, 
            Open_13, Open_14, Open_15, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[19] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[18] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[17] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[16] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[15] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[14] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[13] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[12] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[11] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[10] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[9] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[8] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[7] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[6] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[5] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[4] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[3] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[2] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[1] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi01[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(33)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_5 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, n1142, n1143, n1145, n1147, 
            n1149, n1151, n1153, n1155, n1157, n1159, n1161, n1721}), 
            .B({10'b0000000000, \u_scaler_gray/tdata10[7] , \u_scaler_gray/tdata10[6] , 
            \u_scaler_gray/tdata10[5] , \u_scaler_gray/tdata10[4] , \u_scaler_gray/tdata10[3] , 
            \u_scaler_gray/tdata10[2] , \u_scaler_gray/tdata10[1] , \u_scaler_gray/tdata10[0] }), 
            .O({Open_16, Open_17, Open_18, Open_19, Open_20, Open_21, 
            Open_22, Open_23, Open_24, Open_25, Open_26, Open_27, 
            Open_28, Open_29, Open_30, Open_31, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[19] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[18] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[17] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[16] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[15] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[14] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[13] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[12] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[11] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[10] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[9] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[8] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[7] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[6] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[5] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[4] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[3] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[2] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[1] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi10[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(34)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_6 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b0), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] }), 
            .B({6'b000000, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0] }), 
            .O({Open_32, Open_33, Open_34, Open_35, Open_36, Open_37, 
            Open_38, Open_39, Open_40, Open_41, Open_42, Open_43, 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[23] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[22] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[21] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[20] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[19] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[18] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[17] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[16] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[15] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[14] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[13] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[12] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi00[11] , 
            Open_44, Open_45, Open_46, Open_47, Open_48, Open_49, 
            Open_50, Open_51, Open_52, Open_53, Open_54})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b0, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b0, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(50)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .A_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTA_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_15 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b0), .RSTA(1'b0), .CEB(1'b1), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[10] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcx_fix[0] }), 
            .B({6'b000000, \u_scaler_gray/u1_bilinear_gray/srcy_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[10] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[8] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[7] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[6] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[5] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[4] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[3] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[2] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[1] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[0] }), .O({Open_55, 
            Open_56, Open_57, Open_58, Open_59, Open_60, Open_61, 
            Open_62, Open_63, Open_64, Open_65, Open_66, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[23] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[22] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[21] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[20] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[19] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[18] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[17] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[16] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[15] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[14] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[13] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[12] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi10[11] , 
            Open_67, Open_68, Open_69, Open_70, Open_71, Open_72, 
            Open_73, Open_74, Open_75, Open_76, Open_77})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b0, B_REG=1'b1, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b0, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b1, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(52)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .A_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .B_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTA_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTB_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_17 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b0), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({18'b000001001100110011}), .B({2'b00, \u_scaler_gray/desty[15] , 
            \u_scaler_gray/desty[14] , \u_scaler_gray/desty[13] , \u_scaler_gray/desty[12] , 
            \u_scaler_gray/desty[11] , \u_scaler_gray/desty[10] , \u_scaler_gray/desty[9] , 
            \u_scaler_gray/desty[8] , \u_scaler_gray/desty[7] , \u_scaler_gray/desty[6] , 
            \u_scaler_gray/desty[5] , \u_scaler_gray/desty[4] , \u_scaler_gray/desty[3] , 
            \u_scaler_gray/desty[2] , \u_scaler_gray/desty[1] , \u_scaler_gray/desty[0] }), 
            .O({Open_78, Open_79, Open_80, Open_81, Open_82, Open_83, 
            Open_84, Open_85, \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[27] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[26] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[25] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[24] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[23] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[22] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[21] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[20] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[19] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[18] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[17] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[16] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[15] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[14] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[13] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[12] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[11] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[10] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[9] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[8] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[7] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[6] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[5] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[4] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[3] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[2] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[1] , 
            \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.init_srcy_location[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b0, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b0, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_srcxy.v(55)
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .A_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTA_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/mult_5_pp_0x0 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, n1199, n1200, n1202, n1204, 
            n1206, n1208, n1210, n1212, n1214, n1216, n1218, n1674}), 
            .B({10'b0000000000, \u_scaler_gray/tdata00[7] , \u_scaler_gray/tdata00[6] , 
            \u_scaler_gray/tdata00[5] , \u_scaler_gray/tdata00[4] , \u_scaler_gray/tdata00[3] , 
            \u_scaler_gray/tdata00[2] , \u_scaler_gray/tdata00[1] , \u_scaler_gray/tdata00[0] }), 
            .O({Open_86, Open_87, Open_88, Open_89, Open_90, Open_91, 
            Open_92, Open_93, Open_94, Open_95, Open_96, Open_97, 
            Open_98, Open_99, Open_100, Open_101, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[19] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[18] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[17] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[16] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[15] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[14] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[13] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[12] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[11] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[10] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[9] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[8] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[7] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[6] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[5] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[4] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[3] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[2] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[1] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi00[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(32)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_4 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b1), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, \u_scaler_gray/u1_bilinear_gray/srcx_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/srcx_fix[10] , \u_scaler_gray/u1_bilinear_gray/srcx_fix[9] , 
            9'b000000000}), .B({6'b000000, \u_scaler_gray/u1_bilinear_gray/srcy_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[10] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[8] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[7] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[6] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[5] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[4] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[3] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[2] , \u_scaler_gray/u1_bilinear_gray/srcy_fix[1] , 
            \u_scaler_gray/u1_bilinear_gray/srcy_fix[0] }), .O({Open_102, 
            Open_103, Open_104, Open_105, Open_106, Open_107, Open_108, 
            Open_109, Open_110, Open_111, Open_112, Open_113, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[23] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[22] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[21] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[20] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[19] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[18] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[17] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[16] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[15] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[14] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[13] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[12] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi11[11] , 
            Open_114, Open_115, Open_116, Open_117, Open_118, Open_119, 
            Open_120, Open_121, Open_122, Open_123, Open_124})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b1, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b1, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(53)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .B_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTB_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_18 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, \u_scaler_gray/u1_bilinear_gray/srcx_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/srcx_fix[10] , \u_scaler_gray/u1_bilinear_gray/srcx_fix[9] , 
            9'b000000000}), .B({6'b000000, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[11] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[10] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[9] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[8] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[7] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[6] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[5] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[4] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[3] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[2] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[1] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/comp_srcy_fix[0] }), 
            .O({Open_125, Open_126, Open_127, Open_128, Open_129, 
            Open_130, Open_131, Open_132, Open_133, Open_134, Open_135, 
            Open_136, \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[23] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[22] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[21] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[20] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[19] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[18] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[17] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[16] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[15] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[14] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[13] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[12] , 
            \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/multi01[11] , 
            Open_137, Open_138, Open_139, Open_140, Open_141, Open_142, 
            Open_143, Open_144, Open_145, Open_146, Open_147})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_weight.v(51)
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u1_cal_bilinear_weight/mult_16 .SR_SYNC_PRIORITY = 1'b1;
    EFX_MULT \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7  (.CLK(\Axi_Clk~O ), 
            .CEA(1'b1), .RSTA(1'b0), .CEB(1'b0), .RSTB(1'b0), .CEO(1'b1), 
            .RSTO(1'b0), .A({6'b000000, n1103, n1104, n1106, n1108, 
            n1110, n1114, n1132, n1134, n1136, n1138, n1140, n1723}), 
            .B({10'b0000000000, \u_scaler_gray/tdata11[7] , \u_scaler_gray/tdata11[6] , 
            \u_scaler_gray/tdata11[5] , \u_scaler_gray/tdata11[4] , \u_scaler_gray/tdata11[3] , 
            \u_scaler_gray/tdata11[2] , \u_scaler_gray/tdata11[1] , \u_scaler_gray/tdata11[0] }), 
            .O({Open_148, Open_149, Open_150, Open_151, Open_152, 
            Open_153, Open_154, Open_155, Open_156, Open_157, Open_158, 
            Open_159, Open_160, Open_161, Open_162, Open_163, \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[19] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[18] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[17] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[16] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[15] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[14] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[13] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[12] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[11] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[10] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[9] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[8] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[7] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[6] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[5] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[4] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[3] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[2] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[1] , 
            \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/multi11[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_MULT, WIDTH=18, EFX_ATTRIBUTE_INSTANCE__IS_STF_MULT_PRE_SYNTHESIZED=TRUE, A_REG=1'b1, B_REG=1'b0, O_REG=1'b1, CLK_POLARITY=1'b1, CEA_POLARITY=1'b1, RSTA_POLARITY=1'b1, RSTA_SYNC=1'b1, RSTA_VALUE=1'b0, CEB_POLARITY=1'b1, RSTB_POLARITY=1'b1, RSTB_SYNC=1'b0, RSTB_VALUE=1'b0, CEO_POLARITY=1'b1, RSTO_POLARITY=1'b1, RSTO_SYNC=1'b1, RSTO_VALUE=1'b0, SR_SYNC_PRIORITY=1'b1 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\Bilinear_interpolation\cal_bilinear_data.v(35)
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .WIDTH = 18;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .A_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .B_REG = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .O_REG = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .CLK_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .CEA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTA_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTA_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTA_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .CEB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTB_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTB_SYNC = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTB_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .CEO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTO_POLARITY = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTO_SYNC = 1'b1;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .RSTO_VALUE = 1'b0;
    defparam \u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/mult_7 .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 LUT__10593 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/wdata_cnt_dly[3] ), 
            .O(n7038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10593.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10594 (.I0(n7038), .I1(\u_axi4_ctrl/wdata_cnt_dly[4] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[5] ), .O(n7039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10594.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10595 (.I0(n7039), .I1(\u_axi4_ctrl/wdata_cnt_dly[6] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[5] ), .I3(DdrCtrl_WREADY_0), 
            .O(n7040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hdff3 */ ;
    defparam LUT__10595.LUTMASK = 16'hdff3;
    EFX_LUT4 LUT__10596 (.I0(\u_axi4_ctrl/state[2] ), .I1(\u_axi4_ctrl/state[1] ), 
            .O(DdrCtrl_BREADY_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10596.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10597 (.I0(\u_axi4_ctrl/state[0] ), .I1(DdrCtrl_BREADY_0), 
            .O(DdrCtrl_WVALID_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10597.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10598 (.I0(n7040), .I1(\u_axi4_ctrl/wdata_cnt_dly[7] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[8] ), .I3(DdrCtrl_WVALID_0), 
            .O(n7041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10598.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10599 (.I0(\u_axi4_ctrl/wdata_cnt_dly[3] ), .I1(n7037), 
            .I2(DdrCtrl_WREADY_0), .I3(n7041), .O(DdrCtrl_WLAST_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__10599.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__10600 (.I0(\u_axi4_ctrl/state[1] ), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(\u_axi4_ctrl/state[2] ), .O(DdrCtrl_RREADY_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10600.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10601 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), .O(n7042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10601.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10602 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .O(n7043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__10602.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__10603 (.I0(n7043), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .O(n7044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2fba */ ;
    defparam LUT__10603.LUTMASK = 16'h2fba;
    EFX_LUT4 LUT__10604 (.I0(n7042), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .I2(n7044), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_ctrl_clk ), 
            .O(cmos_sclk)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff0b */ ;
    defparam LUT__10604.LUTMASK = 16'hff0b;
    EFX_LUT4 LUT__10605 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .O(n7045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h233f */ ;
    defparam LUT__10605.LUTMASK = 16'h233f;
    EFX_LUT4 LUT__10606 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .I1(n7044), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .O(n7046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10606.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10607 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I1(n7045), .I2(n7046), .O(cmos_sdat_OE)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__10607.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__10608 (.I0(\PowerOnResetCnt[4] ), .I1(\PowerOnResetCnt[5] ), 
            .I2(\PowerOnResetCnt[6] ), .I3(\PowerOnResetCnt[7] ), .O(n7047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10608.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10609 (.I0(\PowerOnResetCnt[0] ), .I1(\PowerOnResetCnt[1] ), 
            .I2(\PowerOnResetCnt[2] ), .I3(\PowerOnResetCnt[3] ), .O(n7048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10609.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10610 (.I0(n7047), .I1(n7048), .O(\reduce_nand_9/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10610.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10611 (.I0(\u_scaler_gray/srcy_int[0] ), .I1(\u_scaler_gray/srcy_int[1] ), 
            .I2(\u_scaler_gray/srcy_int[2] ), .I3(\u_scaler_gray/srcy_int[3] ), 
            .O(n7049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10611.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10612 (.I0(n7049), .I1(\u_scaler_gray/srcy_int[4] ), .I2(\u_scaler_gray/srcy_int[5] ), 
            .I3(\u_scaler_gray/srcy_int[6] ), .O(n7050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10612.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10613 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] ), 
            .I1(n7050), .I2(\u_scaler_gray/srcy_int[7] ), .O(n7051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__10613.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__10614 (.I0(n7049), .I1(\u_scaler_gray/srcy_int[4] ), .O(n7052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10614.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10615 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] ), 
            .I1(\u_scaler_gray/srcy_int[6] ), .O(n7053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__10615.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__10616 (.I0(n7053), .I1(n7052), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] ), 
            .I3(\u_scaler_gray/srcy_int[5] ), .O(n7054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be */ ;
    defparam LUT__10616.LUTMASK = 16'he7be;
    EFX_LUT4 LUT__10617 (.I0(n7049), .I1(\u_scaler_gray/srcy_int[4] ), .I2(\u_scaler_gray/srcy_int[5] ), 
            .O(n7055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10617.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10618 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] ), 
            .I1(\u_scaler_gray/srcy_int[5] ), .O(n7056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__10618.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__10619 (.I0(n7056), .I1(n7049), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] ), 
            .I3(\u_scaler_gray/srcy_int[4] ), .O(n7057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdd7 */ ;
    defparam LUT__10619.LUTMASK = 16'hbdd7;
    EFX_LUT4 LUT__10620 (.I0(n7055), .I1(n7053), .I2(n7057), .O(n7058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__10620.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__10621 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] ), .I2(n7058), 
            .I3(n7054), .O(n7059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__10621.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__10622 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] ), 
            .I1(\u_scaler_gray/srcy_int[3] ), .O(n7060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__10622.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__10623 (.I0(\u_scaler_gray/srcy_int[0] ), .I1(\u_scaler_gray/srcy_int[1] ), 
            .O(n7061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10623.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10624 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] ), 
            .I1(n7060), .I2(n7061), .I3(\u_scaler_gray/srcy_int[2] ), 
            .O(n7062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__10624.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__10625 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] ), .I2(\u_scaler_gray/srcy_int[0] ), 
            .I3(\u_scaler_gray/srcy_int[1] ), .O(n7063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f75 */ ;
    defparam LUT__10625.LUTMASK = 16'h1f75;
    EFX_LUT4 LUT__10626 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] ), 
            .I1(\u_scaler_gray/srcy_int[1] ), .I2(\u_scaler_gray/srcy_int[2] ), 
            .O(n7064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b */ ;
    defparam LUT__10626.LUTMASK = 16'h2b2b;
    EFX_LUT4 LUT__10627 (.I0(n7064), .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] ), 
            .I2(\u_scaler_gray/srcy_int[3] ), .I3(n7049), .O(n7065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0071 */ ;
    defparam LUT__10627.LUTMASK = 16'h0071;
    EFX_LUT4 LUT__10628 (.I0(n7063), .I1(n7062), .I2(n7065), .I3(n7054), 
            .O(n7066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__10628.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__10629 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] ), 
            .I1(n7059), .I2(n7066), .I3(n7058), .O(n7067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0dcc */ ;
    defparam LUT__10629.LUTMASK = 16'h0dcc;
    EFX_LUT4 LUT__10630 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] ), 
            .I1(\u_scaler_gray/srcy_int[9] ), .O(n7068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__10630.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__10631 (.I0(n7050), .I1(\u_scaler_gray/srcy_int[7] ), .O(n7069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10631.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10632 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] ), 
            .I1(n7068), .I2(n7069), .I3(\u_scaler_gray/srcy_int[8] ), 
            .O(n7070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__10632.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__10633 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] ), 
            .I1(n7050), .I2(\u_scaler_gray/srcy_int[7] ), .I3(n7070), 
            .O(n7071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d */ ;
    defparam LUT__10633.LUTMASK = 16'h007d;
    EFX_LUT4 LUT__10634 (.I0(n7050), .I1(\u_scaler_gray/srcy_int[7] ), .I2(\u_scaler_gray/srcy_int[8] ), 
            .O(n7072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10634.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10635 (.I0(n7072), .I1(\u_scaler_gray/srcy_int[9] ), .O(n7073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10635.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10636 (.I0(\u_scaler_gray/srcy_int[7] ), .I1(n7050), .I2(\u_scaler_gray/srcy_int[8] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] ), .O(n7074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__10636.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__10637 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] ), 
            .I1(n7074), .I2(n7072), .I3(\u_scaler_gray/srcy_int[9] ), 
            .O(n7075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf2ab */ ;
    defparam LUT__10637.LUTMASK = 16'hf2ab;
    EFX_LUT4 LUT__10638 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] ), 
            .I1(n7073), .I2(\u_scaler_gray/srcy_int[10] ), .I3(n7075), 
            .O(n7076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb00 */ ;
    defparam LUT__10638.LUTMASK = 16'heb00;
    EFX_LUT4 LUT__10639 (.I0(n7067), .I1(n7051), .I2(n7071), .I3(n7076), 
            .O(n7077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__10639.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__10640 (.I0(n7072), .I1(\u_scaler_gray/srcy_int[9] ), .I2(\u_scaler_gray/srcy_int[10] ), 
            .O(n7078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10640.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10641 (.I0(n7078), .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] ), 
            .I2(\u_scaler_gray/srcy_int[11] ), .O(n7079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__10641.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__10642 (.I0(n7073), .I1(\u_scaler_gray/srcy_int[10] ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] ), .O(n7080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__10642.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__10643 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] ), 
            .I1(\u_scaler_gray/srcy_int[12] ), .O(n7081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__10643.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__10644 (.I0(n7078), .I1(\u_scaler_gray/srcy_int[11] ), 
            .I2(n7081), .O(n7082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__10644.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__10645 (.I0(n7080), .I1(n7082), .I2(n7079), .O(n7083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10645.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10646 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] ), 
            .I1(n7081), .I2(n7078), .I3(\u_scaler_gray/srcy_int[11] ), 
            .O(n7084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110 */ ;
    defparam LUT__10646.LUTMASK = 16'h0110;
    EFX_LUT4 LUT__10647 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] ), 
            .I1(\u_scaler_gray/srcy_int[13] ), .O(n7085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__10647.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__10648 (.I0(n7078), .I1(\u_scaler_gray/srcy_int[11] ), 
            .I2(\u_scaler_gray/srcy_int[12] ), .I3(n7085), .O(n7086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__10648.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__10649 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] ), 
            .I1(n7082), .I2(n7084), .I3(n7086), .O(n7087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__10649.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__10650 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] ), 
            .I1(\u_scaler_gray/srcy_int[15] ), .O(n7088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__10650.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__10651 (.I0(\u_scaler_gray/srcy_int[10] ), .I1(\u_scaler_gray/srcy_int[11] ), 
            .I2(\u_scaler_gray/srcy_int[12] ), .I3(\u_scaler_gray/srcy_int[13] ), 
            .O(n7089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10651.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10652 (.I0(n7072), .I1(n7089), .I2(\u_scaler_gray/srcy_int[9] ), 
            .O(n7090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10652.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10653 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] ), 
            .I1(n7088), .I2(n7090), .I3(\u_scaler_gray/srcy_int[14] ), 
            .O(n7091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77b */ ;
    defparam LUT__10653.LUTMASK = 16'he77b;
    EFX_LUT4 LUT__10654 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] ), 
            .I1(n7086), .I2(n7091), .O(n7092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__10654.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__10655 (.I0(n7077), .I1(n7083), .I2(n7087), .I3(n7092), 
            .O(n7093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__10655.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__10656 (.I0(n7090), .I1(\u_scaler_gray/srcy_int[14] ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] ), .O(n7094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__10656.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__10657 (.I0(n7094), .I1(\u_scaler_gray/srcy_int[15] ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] ), .O(n7095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__10657.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__10658 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[5] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[4] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[6] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[7] ), .O(n7096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10658.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10659 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[0] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[1] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[2] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[3] ), .O(n7097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10659.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10660 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[12] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[13] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[14] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[15] ), .O(n7098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10660.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10661 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[8] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[10] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[11] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_cnt[9] ), .O(n7099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10661.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10662 (.I0(n7096), .I1(n7097), .I2(n7098), .I3(n7099), 
            .O(n7100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10662.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10663 (.I0(n7095), .I1(n7093), .I2(n7100), .I3(empty), 
            .O(n197_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__10663.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__10664 (.I0(n2741), .I1(n2743), .I2(n2745), .I3(n2747), 
            .O(n7101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10664.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10665 (.I0(n2749), .I1(n2751), .I2(n2753), .I3(n7101), 
            .O(n7102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10665.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10666 (.I0(n2733), .I1(n2735), .I2(n2737), .I3(n2739), 
            .O(n7103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10666.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10667 (.I0(n721), .I1(n2728), .I2(n2729), .I3(n2731), 
            .O(n7104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10667.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10668 (.I0(n7102), .I1(n7103), .I2(n7104), .O(n7105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10668.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10669 (.I0(empty), .I1(n197_2), .I2(n7105), .I3(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), 
            .O(n2105_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__10669.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__10670 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[1] ), .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[0] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/line_cnt[2] ), .I3(\u_CMOS_Capture_RAW_Gray/line_cnt[3] ), 
            .O(n7106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__10670.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__10671 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[4] ), .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[9] ), 
            .I2(n7106), .I3(\u_CMOS_Capture_RAW_Gray/line_cnt[8] ), .O(n7107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00d4 */ ;
    defparam LUT__10671.LUTMASK = 16'h00d4;
    EFX_LUT4 LUT__10672 (.I0(n7107), .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[5] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/line_cnt[8] ), .I3(\u_CMOS_Capture_RAW_Gray/line_cnt[9] ), 
            .O(n7108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf20d */ ;
    defparam LUT__10672.LUTMASK = 16'hf20d;
    EFX_LUT4 LUT__10673 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[8] ), .I1(\u_CMOS_Capture_RAW_Gray/line_cnt[7] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/line_cnt[6] ), .I3(\u_CMOS_Capture_RAW_Gray/line_cnt[9] ), 
            .O(n7109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4001 */ ;
    defparam LUT__10673.LUTMASK = 16'h4001;
    EFX_LUT4 LUT__10674 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[11] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_href_r[1] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/frame_sync_flag ), .I3(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1] ), 
            .O(n7110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10674.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10675 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[10] ), .I1(n7110), 
            .O(n7111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10675.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10676 (.I0(n7109), .I1(n7108), .I2(\u_CMOS_Capture_RAW_Gray/line_cnt[8] ), 
            .I3(n7111), .O(cmos_frame_href)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d00 */ ;
    defparam LUT__10676.LUTMASK = 16'h3d00;
    EFX_LUT4 LUT__10677 (.I0(cmos_frame_href), .I1(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[2] ), 
            .O(\cmos_frame_Gray[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10677.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10678 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][12] ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][13] ), 
            .O(n7112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6996 */ ;
    defparam LUT__10678.LUTMASK = 16'h6996;
    EFX_LUT4 LUT__10679 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2_q ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] ), 
            .O(n7113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__10679.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__10680 (.I0(n7113), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .O(n7114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__10680.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__10681 (.I0(n7114), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .O(n7115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__10681.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__10682 (.I0(n7115), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .O(n7116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__10682.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__10683 (.I0(n7116), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[2] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/waddr[1] ), .O(n7117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1800 */ ;
    defparam LUT__10683.LUTMASK = 16'h1800;
    EFX_LUT4 LUT__10684 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[1] ), .I1(n7116), 
            .I2(\u_afifo_buf/u_efx_fifo_top/waddr[2] ), .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] ), 
            .O(n7118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4001 */ ;
    defparam LUT__10684.LUTMASK = 16'h4001;
    EFX_LUT4 LUT__10685 (.I0(n7117), .I1(n7118), .I2(\u_afifo_buf/u_efx_fifo_top/waddr[0] ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] ), 
            .O(n7119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3553 */ ;
    defparam LUT__10685.LUTMASK = 16'h3553;
    EFX_LUT4 LUT__10686 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[3] ), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .O(n7120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__10686.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__10687 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[5] ), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .O(n7121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__10687.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__10688 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[7] ), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .O(n7122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__10688.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__10689 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13] ), 
            .O(n7123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__10689.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__10690 (.I0(n7123), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/waddr[11] ), .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] ), 
            .O(n7124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77e */ ;
    defparam LUT__10690.LUTMASK = 16'he77e;
    EFX_LUT4 LUT__10691 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF_frt_2_q ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/waddr[10] ), .I2(\u_afifo_buf/u_efx_fifo_top/waddr[9] ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] ), 
            .O(n7125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he77e */ ;
    defparam LUT__10691.LUTMASK = 16'he77e;
    EFX_LUT4 LUT__10692 (.I0(n7124), .I1(n7125), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[13] ), 
            .O(n7126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110 */ ;
    defparam LUT__10692.LUTMASK = 16'h0110;
    EFX_LUT4 LUT__10693 (.I0(n7113), .I1(n7122), .I2(\u_afifo_buf/u_efx_fifo_top/waddr[8] ), 
            .I3(n7126), .O(n7127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8100 */ ;
    defparam LUT__10693.LUTMASK = 16'h8100;
    EFX_LUT4 LUT__10694 (.I0(n7114), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[6] ), 
            .I2(n7121), .I3(n7127), .O(n7128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4200 */ ;
    defparam LUT__10694.LUTMASK = 16'h4200;
    EFX_LUT4 LUT__10695 (.I0(n7115), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[4] ), 
            .I2(n7120), .I3(n7128), .O(n7129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4200 */ ;
    defparam LUT__10695.LUTMASK = 16'h4200;
    EFX_LUT4 LUT__10696 (.I0(n7129), .I1(n7119), .I2(cmos_frame_href), 
            .O(\u_afifo_buf/u_efx_fifo_top/wr_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__10696.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__10697 (.I0(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10697.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10698 (.I0(\r_hdmi_tx0_o[5] ), .I1(\w_hdmi_txd0[0] ), 
            .I2(rc_hdmi_tx), .O(n592_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__10698.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__10699 (.I0(\r_hdmi_tx1_o[5] ), .I1(\w_hdmi_txd1[0] ), 
            .I2(rc_hdmi_tx), .O(n603_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__10699.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__10700 (.I0(\r_hdmi_tx2_o[5] ), .I1(\w_hdmi_txd2[0] ), 
            .I2(rc_hdmi_tx), .O(n614_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__10700.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__10701 (.I0(PllLocked[1]), .I1(PllLocked[0]), .O(n9_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10701.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10702 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] ), .O(n7130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10702.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10703 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] ), .O(n7131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10703.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10704 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] ), .O(n7132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10704.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10705 (.I0(n7130), .I1(n7131), .I2(n7132), .O(n7133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10705.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10706 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] ), .O(n7134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10706.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10707 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] ), .O(n7135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10707.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10708 (.I0(n7133), .I1(n7134), .I2(n7135), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f7f */ ;
    defparam LUT__10708.LUTMASK = 16'h7f7f;
    EFX_LUT4 LUT__10709 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/equal_21/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__10709.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__10710 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__10710.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__10711 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__10711.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10712 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1] ), .O(n7136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10712.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10713 (.I0(n7136), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] ), .O(n7137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10713.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10714 (.I0(n7137), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] ), 
            .O(n7138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__10714.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__10715 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), 
            .I1(n7138), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), 
            .O(n7139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__10715.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__10716 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] ), .O(n7140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10716.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10717 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[3] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[4] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[5] ), .O(n7141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10717.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10718 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[0] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15] ), .O(n7142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10718.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10719 (.I0(n7141), .I1(n7142), .O(n7143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10719.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10720 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[12] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[13] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[14] ), 
            .O(n7144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10720.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10721 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[6] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[7] ), .I2(n7144), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16] ), .O(n7145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10721.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10722 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[8] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[9] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[10] ), 
            .O(n7146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10722.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10723 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[17] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[18] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[19] ), 
            .O(n7147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10723.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10724 (.I0(n7143), .I1(n7145), .I2(n7146), .I3(n7147), 
            .O(n7148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10724.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10725 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[15] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[14] ), .I2(n7148), 
            .O(n7149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10725.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10726 (.I0(n7139), .I1(n7140), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13] ), 
            .I3(n7149), .O(n7150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__10726.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__10727 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] ), 
            .I1(n7150), .O(\u_i2c_timing_ctrl_16reg_16bit/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10727.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10728 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3] ), .O(n7151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10728.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10729 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .O(n7152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10729.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10730 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .O(n7153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10730.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10731 (.I0(n7151), .I1(n7152), .I2(n7153), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .O(n7154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__10731.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__10732 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), .I2(n7151), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .O(n7155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__10732.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__10733 (.I0(n7153), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .O(n7156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10733.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10734 (.I0(n7152), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I2(n7155), .I3(n7156), .O(n7157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__10734.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__10735 (.I0(n7154), .I1(n7157), .O(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10735.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10736 (.I0(n7151), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), .I3(n7153), 
            .O(n7158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__10736.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__10737 (.I0(n7158), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .O(n7159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10737.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10738 (.I0(n7151), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .O(n7160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__10738.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__10739 (.I0(n7151), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .O(n7161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1ff0 */ ;
    defparam LUT__10739.LUTMASK = 16'h1ff0;
    EFX_LUT4 LUT__10740 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), .I2(n7161), 
            .I3(n7152), .O(n7162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__10740.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__10741 (.I0(\i2c_config_index[5] ), .I1(\i2c_config_index[6] ), 
            .I2(\i2c_config_index[7] ), .O(n7163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10741.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10742 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[3] ), 
            .I2(n7163), .O(n7164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__10742.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__10743 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), 
            .O(n7165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10743.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10744 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), .I2(n7164), 
            .I3(n7165), .O(n7166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10744.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10745 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I3(n7151), .O(n7167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbe00 */ ;
    defparam LUT__10745.LUTMASK = 16'hbe00;
    EFX_LUT4 LUT__10746 (.I0(n7167), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), .O(n7168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__10746.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__10747 (.I0(n7148), .I1(n7166), .I2(n7168), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .O(n7169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__10747.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__10748 (.I0(n7160), .I1(n7159), .I2(n7162), .I3(n7169), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__10748.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__10749 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[4] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[3] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[2] ), .O(n7170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10749.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10750 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[1] ), 
            .I1(n7170), .O(n7171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10750.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10751 (.I0(n7171), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), 
            .O(n7172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__10751.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__10752 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), 
            .O(n7173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10752.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10753 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] ), .O(n7174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10753.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10754 (.I0(n7171), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] ), 
            .I2(n7174), .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), 
            .O(n7175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__10754.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__10755 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[13] ), 
            .I1(n7149), .O(n7176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10755.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10756 (.I0(n7175), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] ), .I3(n7176), 
            .O(n7177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7c00 */ ;
    defparam LUT__10756.LUTMASK = 16'h7c00;
    EFX_LUT4 LUT__10757 (.I0(n7172), .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] ), 
            .I2(n7173), .I3(n7177), .O(\u_i2c_timing_ctrl_16reg_16bit/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__10757.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__10758 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[5] ), .I2(n7171), 
            .I3(n7174), .O(n7178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10758.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10759 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), .I2(n7176), 
            .I3(n7178), .O(\u_i2c_timing_ctrl_16reg_16bit/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10759.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10760 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[8] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[9] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[12] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[7] ), .O(n7179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10760.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10761 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[6] ), 
            .I1(n7179), .I2(n7137), .O(n7180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10761.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10762 (.I0(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[11] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/clk_cnt[10] ), .I2(n7176), 
            .I3(n7180), .O(\u_i2c_timing_ctrl_16reg_16bit/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__10762.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__10763 (.I0(\i2c_config_index[0] ), .I1(n7164), .O(\u_i2c_timing_ctrl_16reg_16bit/n205 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10763.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10764 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), .O(n7181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10764.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10765 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), 
            .O(n7182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10765.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10766 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .I2(n7181), 
            .I3(n7182), .O(\u_i2c_timing_ctrl_16reg_16bit/n846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__10766.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__10767 (.I0(n7150), .I1(n3295), .O(\u_i2c_timing_ctrl_16reg_16bit/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10767.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10768 (.I0(n7150), .I1(n3296), .O(\u_i2c_timing_ctrl_16reg_16bit/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10768.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10769 (.I0(n7150), .I1(n3298), .O(\u_i2c_timing_ctrl_16reg_16bit/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10769.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10770 (.I0(n7150), .I1(n3309), .O(\u_i2c_timing_ctrl_16reg_16bit/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10770.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10771 (.I0(n7150), .I1(n3311), .O(\u_i2c_timing_ctrl_16reg_16bit/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10771.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10772 (.I0(n7150), .I1(n3313), .O(\u_i2c_timing_ctrl_16reg_16bit/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10772.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10773 (.I0(n7150), .I1(n3315), .O(\u_i2c_timing_ctrl_16reg_16bit/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10773.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10774 (.I0(n7150), .I1(n3321), .O(\u_i2c_timing_ctrl_16reg_16bit/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10774.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10775 (.I0(n7150), .I1(n3323), .O(\u_i2c_timing_ctrl_16reg_16bit/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10775.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10776 (.I0(n7150), .I1(n3325), .O(\u_i2c_timing_ctrl_16reg_16bit/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10776.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10777 (.I0(n7150), .I1(n3327), .O(\u_i2c_timing_ctrl_16reg_16bit/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10777.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10778 (.I0(n7150), .I1(n3329), .O(\u_i2c_timing_ctrl_16reg_16bit/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10778.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10779 (.I0(n7150), .I1(n3333), .O(\u_i2c_timing_ctrl_16reg_16bit/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10779.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10780 (.I0(n7150), .I1(n3338), .O(\u_i2c_timing_ctrl_16reg_16bit/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10780.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10781 (.I0(n7150), .I1(n219), .O(\u_i2c_timing_ctrl_16reg_16bit/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10781.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10782 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[4] ), .O(n7183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10782.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10783 (.I0(\i2c_config_index[3] ), .I1(n7165), .I2(n7183), 
            .I3(n7163), .O(n7184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10783.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10784 (.I0(n7184), .I1(n7148), .I2(n7156), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .O(n7185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__10784.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__10785 (.I0(n7156), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .O(n7186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10785.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10786 (.I0(n7186), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .O(n7187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__10786.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__10787 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I1(n7156), .I2(n7151), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .O(n7188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfc4 */ ;
    defparam LUT__10787.LUTMASK = 16'hbfc4;
    EFX_LUT4 LUT__10788 (.I0(n7153), .I1(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I2(n7181), .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .O(n7189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__10788.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__10789 (.I0(n7188), .I1(n7189), .O(n7190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10789.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10790 (.I0(n7165), .I1(n7156), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .O(n7191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__10790.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__10791 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .I1(n7191), .O(n7192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10791.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10792 (.I0(n7187), .I1(n7185), .I2(n7190), .I3(n7192), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2 */ ;
    defparam LUT__10792.LUTMASK = 16'hfff2;
    EFX_LUT4 LUT__10793 (.I0(n7148), .I1(n7184), .O(n7193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10793.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10794 (.I0(n7181), .I1(n7191), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), 
            .O(n7194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__10794.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__10795 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I1(n7193), .I2(n7187), .I3(n7194), .O(n7195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__10795.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__10796 (.I0(n7151), .I1(n7186), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[3] ), 
            .I3(n7189), .O(n7196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__10796.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__10797 (.I0(n7195), .I1(n7196), .O(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__10797.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__10798 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n7197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__10798.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__10799 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .O(n7198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10799.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10800 (.I0(n7181), .I1(n7153), .I2(\u_i2c_timing_ctrl_16reg_16bit/current_state[1] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/current_state[4] ), .O(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5780 */ ;
    defparam LUT__10800.LUTMASK = 16'h5780;
    EFX_LUT4 LUT__10801 (.I0(n7197), .I1(n7198), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), .O(n7199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3fa */ ;
    defparam LUT__10801.LUTMASK = 16'hc3fa;
    EFX_LUT4 LUT__10802 (.I0(n7199), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10802.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10803 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), .O(n7200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h32f3 */ ;
    defparam LUT__10803.LUTMASK = 16'h32f3;
    EFX_LUT4 LUT__10804 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I1(n7200), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), 
            .O(ceg_net552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__10804.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__10805 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .O(n7201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdbd */ ;
    defparam LUT__10805.LUTMASK = 16'hbdbd;
    EFX_LUT4 LUT__10806 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(n7201), .O(n7202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10806.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10807 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[2] ), .O(n7203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7fe */ ;
    defparam LUT__10807.LUTMASK = 16'he7fe;
    EFX_LUT4 LUT__10808 (.I0(n7203), .I1(\i2c_config_index[1] ), .O(n7204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10808.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10809 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[1] ), 
            .O(n7205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10809.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10810 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[2] ), 
            .I2(n7205), .I3(\i2c_config_index[4] ), .O(n7206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10810.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10811 (.I0(n7206), .I1(n7204), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I3(n7163), .O(n7207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__10811.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__10812 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(n7206), .I2(n7163), .O(n7208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10812.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10813 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0] ), 
            .I1(n7208), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .O(n7209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__10813.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__10814 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[2] ), .O(n7210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hdcab */ ;
    defparam LUT__10814.LUTMASK = 16'hdcab;
    EFX_LUT4 LUT__10815 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[4] ), .O(n7211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__10815.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__10816 (.I0(n7211), .I1(\i2c_config_index[0] ), .I2(\i2c_config_index[2] ), 
            .O(n7212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10816.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10817 (.I0(n7210), .I1(\i2c_config_index[1] ), .I2(n7212), 
            .I3(n7163), .O(n7213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__10817.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__10818 (.I0(n7213), .I1(n7209), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .O(n7214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__10818.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__10819 (.I0(n7207), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I2(n7214), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n7215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77 */ ;
    defparam LUT__10819.LUTMASK = 16'h0f77;
    EFX_LUT4 LUT__10820 (.I0(n7202), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0] ), 
            .I2(n7215), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h440f */ ;
    defparam LUT__10820.LUTMASK = 16'h440f;
    EFX_LUT4 LUT__10821 (.I0(n7187), .I1(n7185), .I2(n7192), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(n7216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__10821.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__10822 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .I1(n7195), .I2(n7216), .O(n7217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__10822.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__10823 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(n7198), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .O(n7218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__10823.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__10824 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), .O(n7219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10824.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10825 (.I0(n7218), .I1(n7219), .I2(n7217), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), 
            .O(ceg_net664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__10825.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__10826 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .O(n7220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10826.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10827 (.I0(cmos_sdat_IN), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n7221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffc */ ;
    defparam LUT__10827.LUTMASK = 16'h7ffc;
    EFX_LUT4 LUT__10828 (.I0(n7221), .I1(n7220), .I2(n7216), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack5 ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n567 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f50 */ ;
    defparam LUT__10828.LUTMASK = 16'h7f50;
    EFX_LUT4 LUT__10829 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), .O(n7222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10829.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10830 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(n7195), .I2(n7222), .O(n7223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10830.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10831 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .I1(n7223), .O(n7224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10831.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10832 (.I0(n7196), .I1(n7195), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I3(n7222), .O(n7225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__10832.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__10833 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack4 ), .I1(cmos_sdat_IN), 
            .I2(n7224), .I3(n7225), .O(\u_i2c_timing_ctrl_16reg_16bit/n570 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcfa */ ;
    defparam LUT__10833.LUTMASK = 16'hfcfa;
    EFX_LUT4 LUT__10834 (.I0(n7185), .I1(n7187), .O(n7226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10834.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10835 (.I0(n7190), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(n7227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10835.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10836 (.I0(n7227), .I1(n7226), .I2(n7219), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .O(n7228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__10836.LUTMASK = 16'he000;
    EFX_LUT4 LUT__10837 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack3 ), .I1(cmos_sdat_IN), 
            .I2(n7224), .I3(n7228), .O(\u_i2c_timing_ctrl_16reg_16bit/n573 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcfa */ ;
    defparam LUT__10837.LUTMASK = 16'hfcfa;
    EFX_LUT4 LUT__10838 (.I0(n7227), .I1(n7226), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I3(n7219), .O(n7229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__10838.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__10839 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack2 ), .I1(cmos_sdat_IN), 
            .I2(n7224), .I3(n7229), .O(\u_i2c_timing_ctrl_16reg_16bit/n576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcfa */ ;
    defparam LUT__10839.LUTMASK = 16'hfcfa;
    EFX_LUT4 LUT__10840 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I3(n7169), .O(n7230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__10840.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__10841 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack1 ), .I1(cmos_sdat_IN), 
            .I2(n7224), .I3(n7230), .O(\u_i2c_timing_ctrl_16reg_16bit/n579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfcfa */ ;
    defparam LUT__10841.LUTMASK = 16'hfcfa;
    EFX_LUT4 LUT__10842 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), .I2(n7195), 
            .O(n7231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10842.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10843 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack4 ), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack3 ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack2 ), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack1 ), 
            .O(n7232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10843.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10844 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack5 ), .I1(n7231), 
            .I2(n7232), .O(n7233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__10844.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__10845 (.I0(n7162), .I1(n7231), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .O(n7234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__10845.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__10846 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_ack ), .I1(n7233), 
            .I2(n7224), .I3(n7234), .O(\u_i2c_timing_ctrl_16reg_16bit/n581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf3fa */ ;
    defparam LUT__10846.LUTMASK = 16'hf3fa;
    EFX_LUT4 LUT__10847 (.I0(n7146), .I1(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[11] ), 
            .I2(n7144), .I3(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[15] ), 
            .O(n7235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__10847.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__10848 (.I0(\u_i2c_timing_ctrl_16reg_16bit/delay_cnt[16] ), 
            .I1(n7235), .I2(n7147), .O(\u_i2c_timing_ctrl_16reg_16bit/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__10848.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__10849 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), .O(n7236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__10849.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__10850 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .O(n7237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__10850.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__10851 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .O(n7238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf */ ;
    defparam LUT__10851.LUTMASK = 16'ha0cf;
    EFX_LUT4 LUT__10852 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I3(n7238), .O(n7239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a */ ;
    defparam LUT__10852.LUTMASK = 16'hfc0a;
    EFX_LUT4 LUT__10853 (.I0(n7237), .I1(n7236), .I2(n7239), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] ), 
            .O(n7240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10853.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10854 (.I0(n7240), .I1(n7197), .I2(cmos_sdat_OUT), .I3(n7220), 
            .O(n7241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10854.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10855 (.I0(n7240), .I1(cmos_sdat_OUT), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), .O(n7242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc05 */ ;
    defparam LUT__10855.LUTMASK = 16'hfc05;
    EFX_LUT4 LUT__10856 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3] ), .O(n7243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__10856.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__10857 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), .I2(n7240), 
            .I3(n7243), .O(n7244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__10857.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__10858 (.I0(cmos_sdat_OUT), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .O(n7245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h57c5 */ ;
    defparam LUT__10858.LUTMASK = 16'h57c5;
    EFX_LUT4 LUT__10859 (.I0(n7244), .I1(n7242), .I2(n7245), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n7246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__10859.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__10860 (.I0(n7223), .I1(n7241), .I2(n7246), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__10860.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__10861 (.I0(n7169), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I2(n7222), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_transfer_en ), 
            .O(ceg_net632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7d00 */ ;
    defparam LUT__10861.LUTMASK = 16'h7d00;
    EFX_LUT4 LUT__10862 (.I0(n7164), .I1(n222), .O(\u_i2c_timing_ctrl_16reg_16bit/n204 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10862.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10863 (.I0(n7164), .I1(n3293), .O(\u_i2c_timing_ctrl_16reg_16bit/n203 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10863.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10864 (.I0(n3291), .I1(n7164), .O(\u_i2c_timing_ctrl_16reg_16bit/n202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__10864.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__10865 (.I0(n3289), .I1(n7164), .O(\u_i2c_timing_ctrl_16reg_16bit/n201 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__10865.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__10866 (.I0(n7164), .I1(n3287), .O(\u_i2c_timing_ctrl_16reg_16bit/n200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10866.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10867 (.I0(n7164), .I1(n3285), .O(\u_i2c_timing_ctrl_16reg_16bit/n199 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10867.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10868 (.I0(n7164), .I1(n3284), .O(\u_i2c_timing_ctrl_16reg_16bit/n198 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10868.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10869 (.I0(n7199), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .O(\u_i2c_timing_ctrl_16reg_16bit/n499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__10869.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__10870 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .I2(n7199), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] ), .O(\u_i2c_timing_ctrl_16reg_16bit/n498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__10870.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__10871 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[1] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[2] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_stream_cnt[3] ), .O(n7247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__10871.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__10872 (.I0(n7199), .I1(n7247), .O(\u_i2c_timing_ctrl_16reg_16bit/n497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10872.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10873 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[0] ), .O(n7248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc17 */ ;
    defparam LUT__10873.LUTMASK = 16'hfc17;
    EFX_LUT4 LUT__10874 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[4] ), .O(n7249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4ccf */ ;
    defparam LUT__10874.LUTMASK = 16'h4ccf;
    EFX_LUT4 LUT__10875 (.I0(\i2c_config_index[3] ), .I1(n7249), .I2(n7248), 
            .I3(\i2c_config_index[4] ), .O(n7250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heee0 */ ;
    defparam LUT__10875.LUTMASK = 16'heee0;
    EFX_LUT4 LUT__10876 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(n7250), .I2(n7163), .O(n7251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10876.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10877 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[4] ), .O(n7252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb4f */ ;
    defparam LUT__10877.LUTMASK = 16'hfb4f;
    EFX_LUT4 LUT__10878 (.I0(n7252), .I1(n7163), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I3(\i2c_config_index[2] ), .O(n7253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10878.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10879 (.I0(n7253), .I1(n7251), .I2(n7226), .O(n7254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__10879.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__10880 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] ), 
            .I1(n7251), .I2(n7202), .I3(n7217), .O(n7255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__10880.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__10881 (.I0(\i2c_config_index[3] ), .I1(n7205), .I2(\i2c_config_index[2] ), 
            .I3(n7164), .O(n7256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__10881.LUTMASK = 16'he000;
    EFX_LUT4 LUT__10882 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[1] ), .I2(n7256), 
            .I3(n7217), .O(n7257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10882.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10883 (.I0(n7255), .I1(n7254), .I2(n7257), .I3(n7195), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10883.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10884 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[0] ), .O(n7258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ffa */ ;
    defparam LUT__10884.LUTMASK = 16'h3ffa;
    EFX_LUT4 LUT__10885 (.I0(n7258), .I1(\i2c_config_index[4] ), .I2(n7163), 
            .O(n7259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10885.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10886 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[4] ), .I3(\i2c_config_index[2] ), .O(n7260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1700 */ ;
    defparam LUT__10886.LUTMASK = 16'h1700;
    EFX_LUT4 LUT__10887 (.I0(n7252), .I1(n7260), .I2(\i2c_config_index[0] ), 
            .I3(n7163), .O(n7261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1c00 */ ;
    defparam LUT__10887.LUTMASK = 16'h1c00;
    EFX_LUT4 LUT__10888 (.I0(n7261), .I1(n7259), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I3(n7226), .O(n7262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__10888.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__10889 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(n7222), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I3(n7261), .O(n7263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10889.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10890 (.I0(n7202), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] ), 
            .I2(n7263), .I3(n7217), .O(n7264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__10890.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__10891 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[0] ), .O(n7265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10891.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10892 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[2] ), .O(n7266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3001 */ ;
    defparam LUT__10892.LUTMASK = 16'h3001;
    EFX_LUT4 LUT__10893 (.I0(n7266), .I1(n7265), .I2(\i2c_config_index[1] ), 
            .I3(n7163), .O(n7267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__10893.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__10894 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[2] ), .I2(n7267), 
            .I3(n7217), .O(n7268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10894.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10895 (.I0(n7264), .I1(n7262), .I2(n7268), .I3(n7195), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10895.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10896 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[3] ), .O(n7269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3207 */ ;
    defparam LUT__10896.LUTMASK = 16'h3207;
    EFX_LUT4 LUT__10897 (.I0(\i2c_config_index[2] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[1] ), .O(n7270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__10897.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__10898 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[0] ), 
            .I2(n7270), .O(n7271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10898.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10899 (.I0(\i2c_config_index[2] ), .I1(n7269), .I2(n7271), 
            .I3(n7163), .O(n7272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__10899.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__10900 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I1(n7222), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .O(n7273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10900.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10901 (.I0(n7272), .I1(n7273), .I2(n7202), .I3(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3] ), 
            .O(n7274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__10901.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__10902 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .O(n7275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10902.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10903 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[2] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[3] ), .O(n7276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfa3f */ ;
    defparam LUT__10903.LUTMASK = 16'hfa3f;
    EFX_LUT4 LUT__10904 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .O(n7277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10904.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10905 (.I0(\i2c_config_index[3] ), .I1(n7277), .I2(\i2c_config_index[4] ), 
            .I3(\i2c_config_index[0] ), .O(n7278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__10905.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__10906 (.I0(n7276), .I1(\i2c_config_index[1] ), .I2(n7278), 
            .I3(n7163), .O(n7279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__10906.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__10907 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[3] ), .I2(n7279), 
            .I3(n7216), .O(n7280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__10907.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__10908 (.I0(n7275), .I1(n7272), .I2(n7280), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n7281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf077 */ ;
    defparam LUT__10908.LUTMASK = 16'hf077;
    EFX_LUT4 LUT__10909 (.I0(n7281), .I1(n7274), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__10909.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__10910 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[0] ), .I3(\i2c_config_index[1] ), .O(n7282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe3f */ ;
    defparam LUT__10910.LUTMASK = 16'hfe3f;
    EFX_LUT4 LUT__10911 (.I0(\i2c_config_index[2] ), .I1(n7282), .I2(n7164), 
            .O(n7283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__10911.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__10912 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(n7283), .O(n7284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10912.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10913 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I1(n7284), .O(n7285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10913.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10914 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[4] ), 
            .I2(\i2c_config_index[3] ), .O(n7286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3 */ ;
    defparam LUT__10914.LUTMASK = 16'he3e3;
    EFX_LUT4 LUT__10915 (.I0(\i2c_config_index[4] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[3] ), .I3(\i2c_config_index[2] ), .O(n7287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haff3 */ ;
    defparam LUT__10915.LUTMASK = 16'haff3;
    EFX_LUT4 LUT__10916 (.I0(n7286), .I1(\i2c_config_index[1] ), .I2(\i2c_config_index[0] ), 
            .I3(n7287), .O(n7288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10916.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10917 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[4] ), .O(n7289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd08c */ ;
    defparam LUT__10917.LUTMASK = 16'hd08c;
    EFX_LUT4 LUT__10918 (.I0(n7289), .I1(n7183), .I2(\i2c_config_index[3] ), 
            .I3(n7163), .O(n7290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__10918.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__10919 (.I0(n7284), .I1(n7288), .I2(n7290), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .O(n7291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__10919.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__10920 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[4] ), 
            .O(n7292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10920.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10921 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[2] ), 
            .I2(n7292), .I3(n7288), .O(n7293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__10921.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__10922 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4] ), 
            .I1(n7284), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .O(n7294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__10922.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__10923 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), 
            .I1(n7293), .I2(n7163), .I3(n7294), .O(n7295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__10923.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__10924 (.I0(n7291), .I1(n7285), .I2(n7295), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n7296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__10924.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__10925 (.I0(\u_i2c_timing_ctrl_16reg_16bit/current_state[2] ), 
            .I1(n7290), .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[4] ), 
            .I3(n7202), .O(n7297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10925.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10926 (.I0(n7297), .I1(n7296), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__10926.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__10927 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .O(n7298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__10927.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__10928 (.I0(n7205), .I1(n7286), .I2(n7292), .I3(\i2c_config_index[2] ), 
            .O(n7299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10928.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10929 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I1(n7299), .I2(n7163), .O(n7300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10929.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10930 (.I0(n7300), .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5] ), 
            .I2(n7202), .O(n7301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__10930.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10931 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[3] ), 
            .I2(n7277), .O(n7302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__10931.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__10932 (.I0(\i2c_config_index[3] ), .I1(\i2c_config_index[1] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[0] ), .O(n7303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f75 */ ;
    defparam LUT__10932.LUTMASK = 16'h1f75;
    EFX_LUT4 LUT__10933 (.I0(n7302), .I1(n7303), .I2(\i2c_config_index[4] ), 
            .I3(n7163), .O(n7304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8300 */ ;
    defparam LUT__10933.LUTMASK = 16'h8300;
    EFX_LUT4 LUT__10934 (.I0(n7283), .I1(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I2(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[5] ), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .O(n7305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__10934.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__10935 (.I0(n7305), .I1(n7304), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[2] ), .O(n7306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__10935.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__10936 (.I0(n7201), .I1(n7285), .O(n7307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10936.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10937 (.I0(n7300), .I1(n7306), .I2(n7307), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[3] ), 
            .O(n7308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h330e */ ;
    defparam LUT__10937.LUTMASK = 16'h330e;
    EFX_LUT4 LUT__10938 (.I0(n7301), .I1(n7298), .I2(n7308), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__10938.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__10939 (.I0(\i2c_config_index[0] ), .I1(\i2c_config_index[3] ), 
            .I2(\i2c_config_index[1] ), .I3(\i2c_config_index[2] ), .O(n7309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110 */ ;
    defparam LUT__10939.LUTMASK = 16'h0110;
    EFX_LUT4 LUT__10940 (.I0(n7163), .I1(n7309), .I2(\i2c_config_index[4] ), 
            .O(n7310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__10940.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__10941 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6] ), 
            .I1(n7310), .I2(n7273), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(n7311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3533 */ ;
    defparam LUT__10941.LUTMASK = 16'h3533;
    EFX_LUT4 LUT__10942 (.I0(n7195), .I1(n7275), .I2(n7298), .I3(\u_i2c_timing_ctrl_16reg_16bit/next_state[4] ), 
            .O(n7312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__10942.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__10943 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[4] ), .O(n7313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ff2 */ ;
    defparam LUT__10943.LUTMASK = 16'h3ff2;
    EFX_LUT4 LUT__10944 (.I0(\i2c_config_index[4] ), .I1(n7313), .I2(\i2c_config_index[3] ), 
            .I3(n7163), .O(n7314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4300 */ ;
    defparam LUT__10944.LUTMASK = 16'h4300;
    EFX_LUT4 LUT__10945 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[6] ), .I2(n7314), 
            .I3(n7217), .O(n7315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10945.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10946 (.I0(n7315), .I1(n7195), .I2(n7311), .I3(n7312), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h444f */ ;
    defparam LUT__10946.LUTMASK = 16'h444f;
    EFX_LUT4 LUT__10947 (.I0(n7210), .I1(n7205), .I2(n7163), .I3(\i2c_config_index[4] ), 
            .O(n7316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__10947.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__10948 (.I0(n7286), .I1(\i2c_config_index[1] ), .I2(\i2c_config_index[2] ), 
            .I3(n7163), .O(n7317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__10948.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__10949 (.I0(n7317), .I1(n7316), .I2(\u_i2c_timing_ctrl_16reg_16bit/next_state[1] ), 
            .I3(n7226), .O(n7318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__10949.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__10950 (.I0(n7298), .I1(n7217), .O(n7319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10950.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10951 (.I0(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7] ), 
            .I1(n7317), .I2(n7273), .I3(n7319), .O(n7320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__10951.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__10952 (.I0(\i2c_config_index[1] ), .I1(\i2c_config_index[0] ), 
            .I2(\i2c_config_index[2] ), .I3(\i2c_config_index[3] ), .O(n7321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9ef3 */ ;
    defparam LUT__10952.LUTMASK = 16'h9ef3;
    EFX_LUT4 LUT__10953 (.I0(n7321), .I1(n7265), .I2(\i2c_config_index[4] ), 
            .I3(n7163), .O(n7322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc500 */ ;
    defparam LUT__10953.LUTMASK = 16'hc500;
    EFX_LUT4 LUT__10954 (.I0(\u_i2c_timing_ctrl_16reg_16bit/next_state[0] ), 
            .I1(\u_i2c_timing_ctrl_16reg_16bit/i2c_wdata[7] ), .I2(n7322), 
            .I3(n7217), .O(n7323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__10954.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__10955 (.I0(n7320), .I1(n7318), .I2(n7323), .I3(n7195), 
            .O(\u_i2c_timing_ctrl_16reg_16bit/n502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__10955.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__10956 (.I0(\u_rgb2dvi/enc_2/acc[0] ), .I1(\u_rgb2dvi/enc_2/acc[1] ), 
            .I2(\u_rgb2dvi/enc_2/acc[2] ), .I3(\u_rgb2dvi/enc_2/acc[3] ), 
            .O(n7324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__10956.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__10957 (.I0(n7324), .I1(\u_rgb2dvi/enc_2/acc[4] ), .O(n7325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__10957.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__10958 (.I0(\lcd_data[1] ), .I1(\lcd_data[3] ), .O(n7326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__10958.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__10959 (.I0(n7326), .I1(\lcd_data[5] ), .I2(\lcd_data[7] ), 
            .I3(\u_lcd_driver/n133 ), .O(n6895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9600 */ ;
    defparam LUT__10959.LUTMASK = 16'h9600;
    EFX_LUT4 LUT__10960 (.I0(\lcd_data[0] ), .I1(\lcd_data[1] ), .I2(\lcd_data[2] ), 
            .O(n7327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__10960.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__10961 (.I0(n7327), .I1(\lcd_data[3] ), .I2(\lcd_data[4] ), 
            .I3(\u_lcd_driver/n133 ), .O(n7328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6900 */ ;
    defparam LUT__10961.LUTMASK = 16'h6900;
    EFX_LUT4 LUT__10962 (.I0(n7328), .I1(\lcd_data[6] ), .I2(\lcd_data[5] ), 
            .I3(\u_lcd_driver/n133 ), .O(n7329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1777 */ ;
    defparam LUT__10962.LUTMASK = 16'h1777;
    EFX_LUT4 LUT__10963 (.I0(n7327), .I1(\lcd_data[3] ), .I2(\lcd_data[4] ), 
            .O(n7330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b */ ;
    defparam LUT__10963.LUTMASK = 16'h2b2b;
    EFX_LUT4 LUT__10964 (.I0(\lcd_data[3] ), .I1(\lcd_data[4] ), .I2(\lcd_data[5] ), 
            .I3(\lcd_data[6] ), .O(n7331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9669 */ ;
    defparam LUT__10964.LUTMASK = 16'h9669;
    EFX_LUT4 LUT__10965 (.I0(\lcd_data[1] ), .I1(\lcd_data[2] ), .I2(\lcd_data[7] ), 
            .O(n7332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__10965.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__10966 (.I0(\lcd_data[0] ), .I1(\u_lcd_driver/n133 ), .O(n7333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10966.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10967 (.I0(n7331), .I1(n7332), .I2(n7333), .O(n7334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__10967.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__10968 (.I0(\u_lcd_driver/n133 ), .I1(\lcd_data[7] ), .O(n7335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__10968.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__10969 (.I0(n7327), .I1(n7331), .I2(n7335), .O(n7336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__10969.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__10970 (.I0(\lcd_data[0] ), .I1(\lcd_data[1] ), .I2(\lcd_data[2] ), 
            .I3(\u_lcd_driver/n133 ), .O(n7337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he800 */ ;
    defparam LUT__10970.LUTMASK = 16'he800;
    EFX_LUT4 LUT__10971 (.I0(n7330), .I1(n7334), .I2(n7336), .I3(n7337), 
            .O(n7338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eef */ ;
    defparam LUT__10971.LUTMASK = 16'h8eef;
    EFX_LUT4 LUT__10972 (.I0(n7330), .I1(n7336), .I2(n7337), .I3(n7334), 
            .O(n7339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4fd */ ;
    defparam LUT__10972.LUTMASK = 16'hd4fd;
    EFX_LUT4 LUT__10973 (.I0(n7338), .I1(n7329), .I2(n7339), .O(\u_rgb2dvi/enc_0/n103 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__10973.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__10974 (.I0(n7327), .I1(n7331), .I2(\u_lcd_driver/n133 ), 
            .O(n7340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__10974.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__10975 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25_q ), .I2(\u_lcd_driver/r_lcd_dv~FF_frt_7_q ), 
            .O(n7341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__10975.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__10976 (.I0(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q ), 
            .I1(n7341), .O(n7342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10976.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10977 (.I0(n7327), .I1(\u_lcd_driver/n133 ), .O(n7343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__10977.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__10978 (.I0(\lcd_data[0] ), .I1(\lcd_data[1] ), .I2(\u_lcd_driver/n133 ), 
            .O(n7344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__10978.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__10979 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q ), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_19_q ), .O(n7345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8ee8 */ ;
    defparam LUT__10979.LUTMASK = 16'h8ee8;
    EFX_LUT4 LUT__10980 (.I0(n7327), .I1(\lcd_data[3] ), .I2(\u_lcd_driver/n133 ), 
            .O(n7346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__10980.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__10981 (.I0(n7329), .I1(n7338), .I2(n7339), .I3(n7346), 
            .O(n7347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70 */ ;
    defparam LUT__10981.LUTMASK = 16'h8f70;
    EFX_LUT4 LUT__10982 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18_q ), 
            .I2(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_q ), .O(n7348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__10982.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__10983 (.I0(n7329), .I1(n7338), .I2(n7339), .I3(\lcd_data[5] ), 
            .O(n7349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70 */ ;
    defparam LUT__10983.LUTMASK = 16'h8f70;
    EFX_LUT4 LUT__10984 (.I0(\lcd_data[5] ), .I1(\lcd_data[6] ), .I2(n7326), 
            .O(n7350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__10984.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__10985 (.I0(n7326), .I1(\lcd_data[5] ), .I2(\lcd_data[6] ), 
            .I3(\u_lcd_driver/n133 ), .O(n7351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbe00 */ ;
    defparam LUT__10985.LUTMASK = 16'hbe00;
    EFX_LUT4 LUT__10986 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_23_q ), .I2(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_22_q ), 
            .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_q ), .O(n7352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he01f */ ;
    defparam LUT__10986.LUTMASK = 16'he01f;
    EFX_LUT4 LUT__10987 (.I0(n7342), .I1(n7352), .I2(n7345), .I3(n7348), 
            .O(n7353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eef */ ;
    defparam LUT__10987.LUTMASK = 16'h8eef;
    EFX_LUT4 LUT__10988 (.I0(n352), .I1(n378), .I2(n7325), .I3(n7353), 
            .O(n7354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5335 */ ;
    defparam LUT__10988.LUTMASK = 16'h5335;
    EFX_LUT4 LUT__10989 (.I0(n364), .I1(n357), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .O(n7355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__10989.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__10990 (.I0(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25_q ), .I3(\u_lcd_driver/r_lcd_dv~FF_frt_7_q ), 
            .O(n7356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4114 */ ;
    defparam LUT__10990.LUTMASK = 16'h4114;
    EFX_LUT4 LUT__10991 (.I0(n7356), .I1(n7352), .I2(n7348), .I3(n7345), 
            .O(n7357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb66d */ ;
    defparam LUT__10991.LUTMASK = 16'hb66d;
    EFX_LUT4 LUT__10992 (.I0(\u_rgb2dvi/enc_2/acc[4] ), .I1(n7324), .I2(n7357), 
            .I3(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q ), .O(n7358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__10992.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__10993 (.I0(n7355), .I1(n7354), .I2(n7358), .O(n3881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__10993.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__10994 (.I0(n343), .I1(n353), .I2(n7325), .I3(n7353), 
            .O(n7359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3553 */ ;
    defparam LUT__10994.LUTMASK = 16'h3553;
    EFX_LUT4 LUT__10995 (.I0(n365), .I1(n358), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .O(n7360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__10995.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__10996 (.I0(n7360), .I1(n7359), .I2(n7358), .O(n3884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__10996.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__10997 (.I0(n355), .I1(n379), .I2(n7325), .I3(n7353), 
            .O(n7361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5335 */ ;
    defparam LUT__10997.LUTMASK = 16'h5335;
    EFX_LUT4 LUT__10998 (.I0(n367), .I1(n360), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .O(n7362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__10998.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__10999 (.I0(n7362), .I1(n7361), .I2(n7358), .O(n3887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__10999.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11000 (.I0(n3039), .I1(n3207), .I2(n7325), .I3(n7353), 
            .O(n7363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3553 */ ;
    defparam LUT__11000.LUTMASK = 16'h3553;
    EFX_LUT4 LUT__11001 (.I0(n369), .I1(n362), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .O(n7364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11001.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11002 (.I0(n7364), .I1(n7363), .I2(n7358), .O(n3890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11002.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11003 (.I0(\u_rgb2dvi/enc_1/acc[0] ), .I1(\u_rgb2dvi/enc_1/acc[1] ), 
            .I2(\u_rgb2dvi/enc_1/acc[2] ), .I3(\u_rgb2dvi/enc_1/acc[3] ), 
            .O(n7365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11003.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11004 (.I0(n7365), .I1(\u_rgb2dvi/enc_1/acc[4] ), .O(n7366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11004.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11005 (.I0(n352), .I1(n378), .I2(n7366), .I3(n7353), 
            .O(n7367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5335 */ ;
    defparam LUT__11005.LUTMASK = 16'h5335;
    EFX_LUT4 LUT__11006 (.I0(\u_rgb2dvi/enc_1/acc[4] ), .I1(n7365), .I2(n7357), 
            .I3(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q ), .O(n7368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbb0 */ ;
    defparam LUT__11006.LUTMASK = 16'hbbb0;
    EFX_LUT4 LUT__11007 (.I0(n7355), .I1(n7367), .I2(n7368), .O(n3895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11007.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11008 (.I0(n343), .I1(n353), .I2(n7366), .I3(n7353), 
            .O(n7369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3553 */ ;
    defparam LUT__11008.LUTMASK = 16'h3553;
    EFX_LUT4 LUT__11009 (.I0(n7360), .I1(n7369), .I2(n7368), .O(n3898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11009.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11010 (.I0(n355), .I1(n379), .I2(n7366), .I3(n7353), 
            .O(n7370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5335 */ ;
    defparam LUT__11010.LUTMASK = 16'h5335;
    EFX_LUT4 LUT__11011 (.I0(n7362), .I1(n7370), .I2(n7368), .O(n3901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11011.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11012 (.I0(n3039), .I1(n3207), .I2(n7366), .I3(n7353), 
            .O(n7371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3553 */ ;
    defparam LUT__11012.LUTMASK = 16'h3553;
    EFX_LUT4 LUT__11013 (.I0(n7364), .I1(n7371), .I2(n7368), .O(n3904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11013.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11014 (.I0(n7356), .I1(n7348), .I2(n7345), .I3(n7352), 
            .O(n7372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he8fe */ ;
    defparam LUT__11014.LUTMASK = 16'he8fe;
    EFX_LUT4 LUT__11015 (.I0(n7356), .I1(n7348), .I2(n7352), .I3(n7345), 
            .O(n3920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6996 */ ;
    defparam LUT__11015.LUTMASK = 16'h6996;
    EFX_LUT4 LUT__11016 (.I0(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q ), 
            .I1(n3920), .O(n7373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11016.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11017 (.I0(n7372), .I1(n7373), .O(n3913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11017.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11018 (.I0(n7352), .I1(n7345), .I2(n7348), .I3(n7356), 
            .O(n3923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11018.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11019 (.I0(n3923), .I1(n7372), .O(n3926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11019.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11020 (.I0(n7373), .I1(n3926), .O(n3916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11020.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11021 (.I0(n3920), .I1(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q ), 
            .O(n3919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11021.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11022 (.I0(\u_rgb2dvi/enc_0/acc[0] ), .I1(\u_rgb2dvi/enc_0/acc[1] ), 
            .I2(\u_rgb2dvi/enc_0/acc[2] ), .I3(\u_rgb2dvi/enc_0/acc[3] ), 
            .O(n7374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11022.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11023 (.I0(n7374), .I1(\u_rgb2dvi/enc_0/acc[4] ), .O(n7375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11023.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11024 (.I0(n352), .I1(n378), .I2(n7375), .I3(n7353), 
            .O(n7376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5335 */ ;
    defparam LUT__11024.LUTMASK = 16'h5335;
    EFX_LUT4 LUT__11025 (.I0(\u_rgb2dvi/enc_0/acc[4] ), .I1(n7374), .O(n7377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11025.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11026 (.I0(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q ), 
            .I1(n7357), .I2(n7377), .O(n7378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__11026.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__11027 (.I0(n7355), .I1(n7376), .I2(n7378), .O(n3932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11027.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11028 (.I0(n343), .I1(n353), .I2(n7375), .I3(n7353), 
            .O(n7379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3553 */ ;
    defparam LUT__11028.LUTMASK = 16'h3553;
    EFX_LUT4 LUT__11029 (.I0(n7360), .I1(n7379), .I2(n7378), .O(n3935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11029.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11030 (.I0(n355), .I1(n379), .I2(n7375), .I3(n7353), 
            .O(n7380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5335 */ ;
    defparam LUT__11030.LUTMASK = 16'h5335;
    EFX_LUT4 LUT__11031 (.I0(n7362), .I1(n7380), .I2(n7378), .O(n3938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11031.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11032 (.I0(n3039), .I1(n3207), .I2(n7375), .I3(n7353), 
            .O(n7381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3553 */ ;
    defparam LUT__11032.LUTMASK = 16'h3553;
    EFX_LUT4 LUT__11033 (.I0(n7364), .I1(n7381), .I2(n7378), .O(n3941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11033.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11041 (.I0(\u_CMOS_Capture_RAW_Gray/line_cnt[0] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), 
            .O(\u_CMOS_Capture_RAW_Gray/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11041.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11042 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_href_r[1] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_href_r[0] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .O(ceg_net152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__11042.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__11048 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] ), 
            .O(\u_CMOS_Capture_RAW_Gray/n160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11048.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11049 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[1] ), 
            .O(n7383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11049.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11050 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] ), 
            .I2(n7383), .O(ceg_net158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__11050.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__11051 (.I0(n7383), .I1(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] ), 
            .I2(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] ), .O(\u_CMOS_Capture_RAW_Gray/n171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11051.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11071 (.I0(n443), .I1(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), 
            .O(\u_CMOS_Capture_RAW_Gray/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11071.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11072 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3226), 
            .O(\u_CMOS_Capture_RAW_Gray/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11072.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11073 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3224), 
            .O(\u_CMOS_Capture_RAW_Gray/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11073.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11074 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3222), 
            .O(\u_CMOS_Capture_RAW_Gray/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11074.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11075 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3220), 
            .O(\u_CMOS_Capture_RAW_Gray/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11075.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11076 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3218), 
            .O(\u_CMOS_Capture_RAW_Gray/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11076.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11077 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3216), 
            .O(\u_CMOS_Capture_RAW_Gray/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11077.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11078 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3214), 
            .O(\u_CMOS_Capture_RAW_Gray/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11078.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11079 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3212), 
            .O(\u_CMOS_Capture_RAW_Gray/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11079.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11080 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3210), 
            .O(\u_CMOS_Capture_RAW_Gray/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11080.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11081 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_vsync_r[0] ), .I1(n3209), 
            .O(\u_CMOS_Capture_RAW_Gray/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11081.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11082 (.I0(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[0] ), .I1(\u_CMOS_Capture_RAW_Gray/cmos_fps_cnt[1] ), 
            .O(\u_CMOS_Capture_RAW_Gray/n159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__11082.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__11118 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n4132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11118.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11119 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n4135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11119.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11120 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n4138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11120.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11146 (.I0(\u_sensor_frame_count/delay_cnt[6] ), .I1(\u_sensor_frame_count/delay_cnt[5] ), 
            .I2(\u_sensor_frame_count/delay_cnt[1] ), .I3(\u_sensor_frame_count/delay_cnt[11] ), 
            .O(n7399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11146.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11147 (.I0(\u_sensor_frame_count/delay_cnt[3] ), .I1(\u_sensor_frame_count/delay_cnt[2] ), 
            .I2(\u_sensor_frame_count/delay_cnt[0] ), .I3(\u_sensor_frame_count/delay_cnt[10] ), 
            .O(n7400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11147.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11148 (.I0(\u_sensor_frame_count/delay_cnt[9] ), .I1(\u_sensor_frame_count/delay_cnt[8] ), 
            .I2(\u_sensor_frame_count/delay_cnt[7] ), .I3(\u_sensor_frame_count/delay_cnt[4] ), 
            .O(n7401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11148.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11149 (.I0(n7400), .I1(n7401), .I2(n7399), .I3(\u_sensor_frame_count/delay_cnt[12] ), 
            .O(n7402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__11149.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__11150 (.I0(\u_sensor_frame_count/delay_cnt[13] ), .I1(n7402), 
            .I2(\u_sensor_frame_count/delay_cnt[14] ), .O(n7403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__11150.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__11151 (.I0(\u_sensor_frame_count/delay_cnt[17] ), .I1(\u_sensor_frame_count/delay_cnt[18] ), 
            .I2(\u_sensor_frame_count/delay_cnt[19] ), .O(n7404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__11151.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__11152 (.I0(n7403), .I1(\u_sensor_frame_count/delay_cnt[15] ), 
            .I2(\u_sensor_frame_count/delay_cnt[16] ), .I3(n7404), .O(n7405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__11152.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__11153 (.I0(n7405), .I1(\u_sensor_frame_count/delay_cnt[20] ), 
            .I2(\u_sensor_frame_count/delay_cnt[21] ), .I3(\u_sensor_frame_count/delay_cnt[22] ), 
            .O(n7406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11153.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11154 (.I0(\u_sensor_frame_count/delay_cnt[23] ), .I1(n7406), 
            .I2(\u_sensor_frame_count/delay_cnt[24] ), .I3(\u_sensor_frame_count/delay_cnt[25] ), 
            .O(n7407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__11154.LUTMASK = 16'he000;
    EFX_LUT4 LUT__11155 (.I0(\u_sensor_frame_count/delay_cnt[26] ), .I1(n7407), 
            .I2(\u_sensor_frame_count/delay_cnt[27] ), .O(n7408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__11155.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__11156 (.I0(n7408), .I1(n3067), .O(\u_sensor_frame_count/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11156.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11157 (.I0(n7408), .I1(n3069), .O(\u_sensor_frame_count/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11157.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11158 (.I0(n7408), .I1(n3071), .O(\u_sensor_frame_count/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11158.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11159 (.I0(n7408), .I1(n3073), .O(\u_sensor_frame_count/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11159.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11160 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n4176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11160.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11161 (.I0(n7408), .I1(n3075), .O(\u_sensor_frame_count/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11161.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11162 (.I0(n7408), .I1(n3077), .O(\u_sensor_frame_count/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11162.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11163 (.I0(n7408), .I1(n575), .O(\u_sensor_frame_count/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11163.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11164 (.I0(\u_sensor_frame_count/delay_cnt[14] ), .I1(\u_sensor_frame_count/delay_cnt[23] ), 
            .I2(\u_sensor_frame_count/delay_cnt[26] ), .I3(\u_sensor_frame_count/delay_cnt[27] ), 
            .O(n7409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11164.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11165 (.I0(\u_sensor_frame_count/delay_cnt[12] ), .I1(n7409), 
            .I2(n7404), .O(n7410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11165.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11166 (.I0(n7407), .I1(n7410), .O(\u_sensor_frame_count/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__11166.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__11167 (.I0(\u_sensor_frame_count/cmos_fps_cnt[0] ), .I1(\u_sensor_frame_count/n110 ), 
            .O(\u_sensor_frame_count/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11167.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11168 (.I0(\u_sensor_frame_count/cmos_vsync_r[1] ), .I1(\u_sensor_frame_count/cmos_vsync_r[0] ), 
            .I2(\u_sensor_frame_count/n110 ), .O(ceg_net200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__11168.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__11169 (.I0(n7408), .I1(n3079), .O(\u_sensor_frame_count/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11169.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11170 (.I0(n7408), .I1(n3081), .O(\u_sensor_frame_count/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11170.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11171 (.I0(n7408), .I1(\u_sensor_frame_count/delay_cnt[0] ), 
            .O(\u_sensor_frame_count/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11171.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11172 (.I0(empty), .I1(n197_2), .I2(n7105), .I3(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), 
            .O(n2091_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__11172.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__11173 (.I0(cmos_frame_href), .I1(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[0] ), 
            .O(\cmos_frame_Gray[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11173.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11174 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), .I1(\u_afifo_buf/u_efx_fifo_top/wr_en_int ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11174.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11175 (.I0(n7408), .I1(n3054), .O(\u_sensor_frame_count/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11175.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11176 (.I0(n7408), .I1(n3052), .O(\u_sensor_frame_count/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11176.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11177 (.I0(n7408), .I1(n3047), .O(\u_sensor_frame_count/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11177.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11178 (.I0(n7408), .I1(n3045), .O(\u_sensor_frame_count/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11178.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11179 (.I0(n7408), .I1(n3041), .O(\u_sensor_frame_count/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11179.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11180 (.I0(n7408), .I1(n3037), .O(\u_sensor_frame_count/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11180.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11181 (.I0(n7408), .I1(n3035), .O(\u_sensor_frame_count/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11181.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11182 (.I0(n7408), .I1(n3031), .O(\u_sensor_frame_count/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11182.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11183 (.I0(n7408), .I1(n2900), .O(\u_sensor_frame_count/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11183.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11184 (.I0(n7408), .I1(n2898), .O(\u_sensor_frame_count/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11184.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11185 (.I0(n7408), .I1(n2881), .O(\u_sensor_frame_count/n55 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11185.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11186 (.I0(n7408), .I1(n2879), .O(\u_sensor_frame_count/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11186.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11187 (.I0(n7408), .I1(n2877), .O(\u_sensor_frame_count/n53 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11187.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11188 (.I0(n7408), .I1(n2875), .O(\u_sensor_frame_count/n52 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11188.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11189 (.I0(n7408), .I1(n2873), .O(\u_sensor_frame_count/n51 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11189.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11190 (.I0(n7408), .I1(n2871), .O(\u_sensor_frame_count/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11190.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11191 (.I0(n7408), .I1(n2869), .O(\u_sensor_frame_count/n49 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11191.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11192 (.I0(n7408), .I1(n2868), .O(\u_sensor_frame_count/n48 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11192.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11193 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n4211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11193.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11194 (.I0(\u_sensor_frame_count/n110 ), .I1(n601), .O(\u_sensor_frame_count/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11194.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11195 (.I0(\u_sensor_frame_count/n110 ), .I1(n2866), .O(\u_sensor_frame_count/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11195.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11196 (.I0(\u_sensor_frame_count/n110 ), .I1(n2864), .O(\u_sensor_frame_count/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11196.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11197 (.I0(\u_sensor_frame_count/n110 ), .I1(n2862), .O(\u_sensor_frame_count/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11197.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11198 (.I0(\u_sensor_frame_count/n110 ), .I1(n2860), .O(\u_sensor_frame_count/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11198.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11199 (.I0(\u_sensor_frame_count/n110 ), .I1(n2858), .O(\u_sensor_frame_count/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11199.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11200 (.I0(\u_sensor_frame_count/n110 ), .I1(n2856), .O(\u_sensor_frame_count/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11200.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11201 (.I0(\u_sensor_frame_count/n110 ), .I1(n2855), .O(\u_sensor_frame_count/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11201.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11202 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n4222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11202.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11203 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n4225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11203.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11204 (.I0(empty), .I1(n197_2), .I2(n7105), .O(\u_afifo_buf/u_efx_fifo_top/rd_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__11204.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__11205 (.I0(cmos_frame_href), .I1(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[1] ), 
            .O(\cmos_frame_Gray[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11205.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11206 (.I0(cmos_frame_href), .I1(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[3] ), 
            .O(\cmos_frame_Gray[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11206.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11207 (.I0(cmos_frame_href), .I1(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[4] ), 
            .O(\cmos_frame_Gray[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11207.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11208 (.I0(cmos_frame_href), .I1(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[5] ), 
            .O(\cmos_frame_Gray[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11208.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11209 (.I0(cmos_frame_href), .I1(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[6] ), 
            .O(\cmos_frame_Gray[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11209.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11210 (.I0(cmos_frame_href), .I1(\u_CMOS_Capture_RAW_Gray/cmos_data_r1[7] ), 
            .O(\cmos_frame_Gray[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11210.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11211 (.I0(empty), .I1(n7105), .I2(n197_2), .O(ceg_net219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__11211.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__11212 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][13] ), 
            .O(n6308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11212.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11213 (.I0(n6308), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11] ), 
            .O(n6311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11213.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11214 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_frt_1_q ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10] ), 
            .O(n6314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11214.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11215 (.I0(n6314), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] ), 
            .O(n6317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11215.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11216 (.I0(n6317), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .O(n6320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11216.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11217 (.I0(n6320), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .O(n6326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__11217.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__11218 (.I0(n6326), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .O(n6332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__11218.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__11219 (.I0(n6332), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] ), 
            .I3(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .O(n6341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6996 */ ;
    defparam LUT__11219.LUTMASK = 16'h6996;
    EFX_LUT4 LUT__11220 (.I0(n6341), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] ), 
            .O(n4296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11220.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11221 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .O(n7411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11221.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11222 (.I0(n7411), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[0] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[1] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11222.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11223 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[0] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[1] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11223.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11226 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .O(n7412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11226.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11227 (.I0(n7412), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[1] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[2] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11227.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11228 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .O(n7413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11228.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11229 (.I0(n7413), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[2] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[3] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11229.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11230 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .O(n7414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11230.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11231 (.I0(n7414), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[3] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[4] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11231.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11232 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .O(n7415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11232.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11233 (.I0(n7415), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[4] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[5] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11233.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11234 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .O(n7416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11234.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11235 (.I0(n7416), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[5] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[6] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11235.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11236 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .O(n7417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11236.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11237 (.I0(n7417), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[6] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[7] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11237.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11238 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .O(n7418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11238.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11239 (.I0(n7418), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[7] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[8] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11239.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11240 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .O(n7419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11240.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11241 (.I0(n7419), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[8] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[9] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11241.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11242 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] ), 
            .O(n7420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11242.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11243 (.I0(n7420), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[9] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[10] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11243.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11244 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] ), 
            .O(n7421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11244.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11245 (.I0(n7421), .I1(\u_afifo_buf/u_efx_fifo_top/raddr[10] ), 
            .I2(\u_afifo_buf/u_efx_fifo_top/raddr[11] ), .I3(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11245.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11246 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/raddr[12] ), .I2(empty), .O(n7422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11246.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11247 (.I0(\u_afifo_buf/u_efx_fifo_top/raddr[11] ), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] ), 
            .I2(empty), .I3(n7422), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53 */ ;
    defparam LUT__11247.LUTMASK = 16'hac53;
    EFX_LUT4 LUT__11248 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[13] ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[13] ), 
            .I2(empty), .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11248.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11249 (.I0(n7422), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[13] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11249.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11250 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[1] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[2] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11250.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11251 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[3] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[2] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11251.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11252 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[4] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[3] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11252.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11253 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[5] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[4] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11253.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11254 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[6] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[5] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11254.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11255 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[7] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[6] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11255.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11256 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[8] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[7] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11256.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11257 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[9] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[8] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11257.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11258 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[9] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[10] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11258.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11259 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[10] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[11] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11259.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11260 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[11] ), .I1(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11260.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11261 (.I0(\u_afifo_buf/u_efx_fifo_top/waddr[12] ), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[13] ), 
            .O(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11261.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11262 (.I0(tvalid_o), .I1(\u_scaler_gray/tvalid_o_r ), 
            .O(ceg_net226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11262.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11263 (.I0(\u_scaler_gray/vs_cnt[12] ), .I1(\u_scaler_gray/vs_cnt[13] ), 
            .I2(\u_scaler_gray/vs_cnt[14] ), .I3(\u_scaler_gray/vs_cnt[15] ), 
            .O(n7423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11263.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11264 (.I0(\u_scaler_gray/vs_cnt[7] ), .I1(\u_scaler_gray/vs_cnt[8] ), 
            .I2(\u_scaler_gray/vs_cnt[10] ), .I3(\u_scaler_gray/vs_cnt[11] ), 
            .O(n7424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11264.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11265 (.I0(\u_scaler_gray/vs_cnt[3] ), .I1(\u_scaler_gray/vs_cnt[5] ), 
            .I2(n7423), .I3(n7424), .O(n7425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11265.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11266 (.I0(\u_scaler_gray/vs_cnt[4] ), .I1(\u_scaler_gray/vs_cnt[6] ), 
            .I2(\u_scaler_gray/vs_cnt[9] ), .I3(tvalid_o), .O(n7426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11266.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11267 (.I0(\u_scaler_gray/vs_cnt[0] ), .I1(\u_scaler_gray/tvalid_o_r ), 
            .I2(\u_scaler_gray/vs_cnt[1] ), .I3(\u_scaler_gray/vs_cnt[2] ), 
            .O(n7427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11267.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11268 (.I0(n7425), .I1(n7426), .I2(n7427), .O(\u_scaler_gray/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11268.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11269 (.I0(\u_scaler_gray/vs_cnt[2] ), .I1(\u_scaler_gray/vs_cnt[4] ), 
            .I2(\u_scaler_gray/vs_cnt[6] ), .I3(\u_scaler_gray/vs_cnt[9] ), 
            .O(n7428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11269.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11270 (.I0(n7428), .I1(\u_scaler_gray/vs_cnt[0] ), .I2(\u_scaler_gray/vs_cnt[1] ), 
            .O(n7429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11270.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11271 (.I0(ceg_net226), .I1(n7429), .I2(n7425), .O(n7430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11271.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11272 (.I0(\u_scaler_gray/n150 ), .I1(n7430), .O(ceg_net229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11272.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11273 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[4] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[5] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[6] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[7] ), .O(n7431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11273.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11274 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[0] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[1] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[2] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[3] ), .O(n7432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11274.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11275 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[12] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[13] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[14] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[15] ), .O(n7433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11275.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11276 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[8] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[9] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[11] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_row_pixel_cnt[10] ), .O(n7434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11276.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11277 (.I0(n7431), .I1(n7432), .I2(n7433), .I3(n7434), 
            .O(n7435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11277.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11278 (.I0(n197_2), .I1(n7435), .O(\u_scaler_gray/u0_data_stream_ctr/w_image_tlast )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11278.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11279 (.I0(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .I3(\Axi0ResetReg[2] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1703 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h80ff */ ;
    defparam LUT__11279.LUTMASK = 16'h80ff;
    EFX_LUT4 LUT__11280 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[4] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_addra[5] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_addra[6] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_addra[7] ), .O(n7436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11280.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11281 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[12] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_addra[13] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_addra[14] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_addra[15] ), .O(n7437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11281.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11282 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[9] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_addra[10] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_addra[0] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_addra[11] ), .O(n7438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11282.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11283 (.I0(\u_scaler_gray/u0_data_stream_ctr/w_addra[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/w_addra[2] ), .I2(\u_scaler_gray/u0_data_stream_ctr/w_addra[3] ), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/w_addra[8] ), .O(n7439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11283.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11284 (.I0(n7436), .I1(n7437), .I2(n7438), .I3(n7439), 
            .O(n7440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11284.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11285 (.I0(n7440), .I1(n197_2), .I2(\Axi0ResetReg[2] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1704 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f */ ;
    defparam LUT__11285.LUTMASK = 16'h8f8f;
    EFX_LUT4 LUT__11286 (.I0(n7100), .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), .I3(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), 
            .O(n7441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he033 */ ;
    defparam LUT__11286.LUTMASK = 16'he033;
    EFX_LUT4 LUT__11287 (.I0(\u_scaler_gray/desty[12] ), .I1(\u_scaler_gray/desty[13] ), 
            .I2(\u_scaler_gray/desty[14] ), .I3(\u_scaler_gray/desty[15] ), 
            .O(n7442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11287.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11288 (.I0(\u_scaler_gray/desty[7] ), .I1(\u_scaler_gray/desty[8] ), 
            .I2(\u_scaler_gray/desty[10] ), .I3(\u_scaler_gray/desty[11] ), 
            .O(n7443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11288.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11289 (.I0(\u_scaler_gray/desty[3] ), .I1(\u_scaler_gray/desty[5] ), 
            .I2(n7442), .I3(n7443), .O(n7444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11289.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11290 (.I0(\u_scaler_gray/desty[2] ), .I1(\u_scaler_gray/desty[4] ), 
            .I2(\u_scaler_gray/desty[6] ), .I3(\u_scaler_gray/desty[9] ), 
            .O(n7445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11290.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11291 (.I0(\u_scaler_gray/desty[0] ), .I1(\u_scaler_gray/desty[1] ), 
            .I2(n7444), .I3(n7445), .O(n7446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11291.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11292 (.I0(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[0] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[1] ), .I2(n7446), 
            .I3(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), .O(n7447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__11292.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__11293 (.I0(\u_scaler_gray/srcy_int[8] ), .I1(\u_scaler_gray/srcy_int[10] ), 
            .I2(\u_scaler_gray/srcy_int[11] ), .I3(\u_scaler_gray/srcy_int[9] ), 
            .O(n7448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11293.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11294 (.I0(\u_scaler_gray/srcy_int[4] ), .I1(\u_scaler_gray/srcy_int[5] ), 
            .I2(\u_scaler_gray/srcy_int[6] ), .I3(\u_scaler_gray/srcy_int[7] ), 
            .O(n7449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11294.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11295 (.I0(\u_scaler_gray/srcy_int[12] ), .I1(\u_scaler_gray/srcy_int[13] ), 
            .I2(\u_scaler_gray/srcy_int[14] ), .I3(\u_scaler_gray/srcy_int[15] ), 
            .O(n7450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11295.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11296 (.I0(n7049), .I1(n7448), .I2(n7449), .I3(n7450), 
            .O(n7451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11296.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11297 (.I0(n7451), .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), 
            .O(n7452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11297.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11298 (.I0(\u_scaler_gray/destx[4] ), .I1(\u_scaler_gray/destx[5] ), 
            .I2(\u_scaler_gray/destx[6] ), .I3(\u_scaler_gray/destx[7] ), 
            .O(n7453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11298.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11299 (.I0(\u_scaler_gray/destx[0] ), .I1(\u_scaler_gray/destx[1] ), 
            .I2(\u_scaler_gray/destx[2] ), .I3(\u_scaler_gray/destx[3] ), 
            .O(n7454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11299.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11300 (.I0(\u_scaler_gray/destx[12] ), .I1(\u_scaler_gray/destx[13] ), 
            .I2(\u_scaler_gray/destx[14] ), .I3(\u_scaler_gray/destx[15] ), 
            .O(n7455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11300.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11301 (.I0(\u_scaler_gray/destx[10] ), .I1(\u_scaler_gray/destx[11] ), 
            .I2(\u_scaler_gray/destx[8] ), .I3(\u_scaler_gray/destx[9] ), 
            .O(n7456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11301.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11302 (.I0(n7453), .I1(n7454), .I2(n7455), .I3(n7456), 
            .O(n7457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11302.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11303 (.I0(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), 
            .I1(n7457), .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .O(n7458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__11303.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__11304 (.I0(n7093), .I1(n7095), .I2(n7452), .I3(n7458), 
            .O(n7459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__11304.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__11305 (.I0(n7459), .I1(n7447), .I2(n7441), .I3(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fae */ ;
    defparam LUT__11305.LUTMASK = 16'h0fae;
    EFX_LUT4 LUT__11306 (.I0(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[0] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), .O(\u_scaler_gray/u0_data_stream_ctr/n2156 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11306.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11307 (.I0(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .I3(\Axi0ResetReg[2] ), .O(ceg_net526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbeaa */ ;
    defparam LUT__11307.LUTMASK = 16'hbeaa;
    EFX_LUT4 LUT__11308 (.I0(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__11308.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__11309 (.I0(\u_scaler_gray/u0_data_stream_ctr/equal_59/n5 ), 
            .I1(n7457), .O(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11309.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11310 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
            .I1(\Axi0ResetReg[2] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11310.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11311 (.I0(\u_scaler_gray/desty[2] ), .I1(\u_scaler_gray/desty[4] ), 
            .I2(\u_scaler_gray/desty[6] ), .I3(\u_scaler_gray/desty[9] ), 
            .O(n7460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11311.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11312 (.I0(n7444), .I1(n7460), .I2(\u_scaler_gray/desty[0] ), 
            .I3(\u_scaler_gray/desty[1] ), .O(n7461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11312.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11313 (.I0(n7461), .I1(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
            .I2(\Axi0ResetReg[2] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1713 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f */ ;
    defparam LUT__11313.LUTMASK = 16'h8f8f;
    EFX_LUT4 LUT__11314 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n87 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n86 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11314.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11315 (.I0(\u_scaler_gray/srcx_int[0] ), .I1(\u_scaler_gray/srcx_int[1] ), 
            .O(n7462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11315.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11316 (.I0(\u_scaler_gray/srcx_int[4] ), .I1(\u_scaler_gray/srcx_int[5] ), 
            .I2(\u_scaler_gray/srcx_int[6] ), .I3(\u_scaler_gray/srcx_int[7] ), 
            .O(n7463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11316.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11317 (.I0(n7462), .I1(n7463), .I2(\u_scaler_gray/srcx_int[2] ), 
            .I3(\u_scaler_gray/srcx_int[3] ), .O(n7464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11317.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11318 (.I0(\u_scaler_gray/srcx_int[12] ), .I1(\u_scaler_gray/srcx_int[13] ), 
            .I2(\u_scaler_gray/srcx_int[14] ), .I3(\u_scaler_gray/srcx_int[15] ), 
            .O(n7465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11318.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11319 (.I0(\u_scaler_gray/srcx_int[8] ), .I1(\u_scaler_gray/srcx_int[9] ), 
            .I2(\u_scaler_gray/srcx_int[11] ), .I3(\u_scaler_gray/srcx_int[10] ), 
            .O(n7466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11319.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11320 (.I0(n7465), .I1(n7466), .O(n7467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11320.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11321 (.I0(n7464), .I1(n7467), .O(n7468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11321.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11322 (.I0(n7468), .I1(\u_scaler_gray/srcx_int[0] ), .O(\u_scaler_gray/u0_data_stream_ctr/n903 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11322.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11323 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n102 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n101 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11323.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11324 (.I0(n7435), .I1(n197_2), .I2(\Axi0ResetReg[2] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1702 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f */ ;
    defparam LUT__11324.LUTMASK = 16'h8f8f;
    EFX_LUT4 LUT__11325 (.I0(n7100), .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), .I3(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .O(n7469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf70 */ ;
    defparam LUT__11325.LUTMASK = 16'hcf70;
    EFX_LUT4 LUT__11326 (.I0(n7447), .I1(\u_scaler_gray/u0_data_stream_ctr/r_image_tlast ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), .I3(n7469), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcefc */ ;
    defparam LUT__11326.LUTMASK = 16'hcefc;
    EFX_LUT4 LUT__11327 (.I0(n7446), .I1(\u_scaler_gray/u0_data_stream_ctr/scaler_st[2] ), 
            .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[0] ), .I3(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ecc */ ;
    defparam LUT__11327.LUTMASK = 16'h0ecc;
    EFX_LUT4 LUT__11328 (.I0(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[0] ), 
            .I1(\u_scaler_gray/u0_data_stream_ctr/delay_cnt[1] ), .I2(\u_scaler_gray/u0_data_stream_ctr/scaler_st[1] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n2073 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__11328.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__11329 (.I0(\u_scaler_gray/srcx_int[8] ), .I1(\u_scaler_gray/srcy_int[0] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1196 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11329.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11330 (.I0(\u_scaler_gray/srcx_int[8] ), .I1(\u_scaler_gray/srcy_int[0] ), 
            .I2(\u_scaler_gray/srcx_int[9] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1161 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11330.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11331 (.I0(\u_scaler_gray/srcx_int[8] ), .I1(\u_scaler_gray/srcx_int[9] ), 
            .O(n7470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11331.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11332 (.I0(n7470), .I1(\u_scaler_gray/srcy_int[0] ), .I2(\u_scaler_gray/srcx_int[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1160 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__11332.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__11333 (.I0(n7470), .I1(\u_scaler_gray/srcx_int[10] ), 
            .I2(\u_scaler_gray/srcy_int[0] ), .I3(\u_scaler_gray/srcx_int[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1159 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1fe0 */ ;
    defparam LUT__11333.LUTMASK = 16'h1fe0;
    EFX_LUT4 LUT__11334 (.I0(\u_scaler_gray/u0_data_stream_ctr/n903 ), .I1(\u_scaler_gray/srcx_int[1] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n885 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11334.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11335 (.I0(n7468), .I1(n7462), .I2(\u_scaler_gray/srcx_int[2] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n884 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__11335.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__11336 (.I0(n7468), .I1(n7462), .I2(\u_scaler_gray/srcx_int[2] ), 
            .I3(\u_scaler_gray/srcx_int[3] ), .O(\u_scaler_gray/u0_data_stream_ctr/n883 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfc0 */ ;
    defparam LUT__11336.LUTMASK = 16'hbfc0;
    EFX_LUT4 LUT__11337 (.I0(n7468), .I1(n7462), .I2(\u_scaler_gray/srcx_int[2] ), 
            .I3(\u_scaler_gray/srcx_int[3] ), .O(n7471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__11337.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__11338 (.I0(n7471), .I1(\u_scaler_gray/srcx_int[4] ), .O(\u_scaler_gray/u0_data_stream_ctr/n882 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11338.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11339 (.I0(n7471), .I1(\u_scaler_gray/srcx_int[4] ), .O(n7472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11339.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11340 (.I0(n7472), .I1(\u_scaler_gray/srcx_int[5] ), .O(\u_scaler_gray/u0_data_stream_ctr/n881 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11340.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11341 (.I0(n7472), .I1(\u_scaler_gray/srcx_int[5] ), .O(n7473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11341.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11342 (.I0(n7473), .I1(\u_scaler_gray/srcx_int[6] ), .O(\u_scaler_gray/u0_data_stream_ctr/n880 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11342.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11343 (.I0(n7473), .I1(\u_scaler_gray/srcx_int[6] ), .I2(\u_scaler_gray/srcx_int[7] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n879 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11343.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11344 (.I0(n7467), .I1(n7464), .O(n7474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11344.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11345 (.I0(n7474), .I1(\u_scaler_gray/u0_data_stream_ctr/n1196 ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11345.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11346 (.I0(n7474), .I1(\u_scaler_gray/srcx_int[8] ), .I2(\u_scaler_gray/srcy_int[0] ), 
            .I3(\u_scaler_gray/srcx_int[9] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h17e8 */ ;
    defparam LUT__11346.LUTMASK = 16'h17e8;
    EFX_LUT4 LUT__11347 (.I0(\u_scaler_gray/srcx_int[9] ), .I1(\u_scaler_gray/srcx_int[8] ), 
            .I2(n7464), .I3(\u_scaler_gray/srcy_int[0] ), .O(n7475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha87f */ ;
    defparam LUT__11347.LUTMASK = 16'ha87f;
    EFX_LUT4 LUT__11348 (.I0(n7475), .I1(\u_scaler_gray/srcx_int[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1177 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11348.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11349 (.I0(\u_scaler_gray/srcy_int[0] ), .I1(\u_scaler_gray/srcx_int[10] ), 
            .I2(n7475), .I3(\u_scaler_gray/srcx_int[11] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1176 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h53ac */ ;
    defparam LUT__11349.LUTMASK = 16'h53ac;
    EFX_LUT4 LUT__11350 (.I0(\u_scaler_gray/srcy_int[0] ), .I1(\u_scaler_gray/srcx_int[8] ), 
            .I2(\u_scaler_gray/srcx_int[9] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1195 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__11350.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__11351 (.I0(n7470), .I1(\u_scaler_gray/srcy_int[0] ), .I2(\u_scaler_gray/srcx_int[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1194 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1e1 */ ;
    defparam LUT__11351.LUTMASK = 16'he1e1;
    EFX_LUT4 LUT__11352 (.I0(n7470), .I1(\u_scaler_gray/srcx_int[10] ), 
            .I2(\u_scaler_gray/srcy_int[0] ), .I3(\u_scaler_gray/srcx_int[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1193 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf10e */ ;
    defparam LUT__11352.LUTMASK = 16'hf10e;
    EFX_LUT4 LUT__11353 (.I0(n7474), .I1(\u_scaler_gray/srcx_int[8] ), .I2(\u_scaler_gray/srcy_int[0] ), 
            .I3(\u_scaler_gray/srcx_int[9] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1212 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h718e */ ;
    defparam LUT__11353.LUTMASK = 16'h718e;
    EFX_LUT4 LUT__11354 (.I0(\u_scaler_gray/srcx_int[9] ), .I1(\u_scaler_gray/srcx_int[8] ), 
            .I2(n7464), .I3(\u_scaler_gray/srcy_int[0] ), .O(n7476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fa8 */ ;
    defparam LUT__11354.LUTMASK = 16'h7fa8;
    EFX_LUT4 LUT__11355 (.I0(n7476), .I1(\u_scaler_gray/srcx_int[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/n1211 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11355.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11356 (.I0(\u_scaler_gray/srcy_int[0] ), .I1(\u_scaler_gray/srcx_int[10] ), 
            .I2(n7476), .I3(\u_scaler_gray/srcx_int[11] ), .O(\u_scaler_gray/u0_data_stream_ctr/n1210 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha35c */ ;
    defparam LUT__11356.LUTMASK = 16'ha35c;
    EFX_LUT4 LUT__11357 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n90 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n89 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11357.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11358 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n84 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n83 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11358.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11359 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n93 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n92 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11359.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11360 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n99 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n98 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11360.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11361 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n96 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n95 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11361.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11362 (.I0(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n104 ), 
            .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n105 ), .I2(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ram/n80 ), 
            .O(\tdata_i[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__11362.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__11363 (.I0(n7430), .I1(n900), .O(\u_scaler_gray/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11363.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11364 (.I0(n7430), .I1(n2582), .O(\u_scaler_gray/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11364.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11365 (.I0(n7430), .I1(n2580), .O(\u_scaler_gray/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11365.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11366 (.I0(n7430), .I1(n2578), .O(\u_scaler_gray/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11366.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11367 (.I0(n7430), .I1(n2576), .O(\u_scaler_gray/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11367.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11368 (.I0(n7430), .I1(n2574), .O(\u_scaler_gray/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11368.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11369 (.I0(n7430), .I1(n2572), .O(\u_scaler_gray/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11369.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11370 (.I0(n7430), .I1(n2570), .O(\u_scaler_gray/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11370.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11371 (.I0(n7430), .I1(n2568), .O(\u_scaler_gray/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11371.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11372 (.I0(n7430), .I1(n2566), .O(\u_scaler_gray/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11372.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11373 (.I0(n7430), .I1(n2564), .O(\u_scaler_gray/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11373.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11374 (.I0(n7430), .I1(n2562), .O(\u_scaler_gray/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11374.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11375 (.I0(n7430), .I1(n2548), .O(\u_scaler_gray/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11375.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11376 (.I0(n7430), .I1(n2546), .O(\u_scaler_gray/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11376.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11377 (.I0(n7430), .I1(n2545), .O(\u_scaler_gray/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11377.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11378 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[16] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[17] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[19] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[27] ), 
            .O(n7477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11378.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11379 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[24] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[25] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[26] ), 
            .I3(n7477), .O(n7478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11379.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11380 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[12] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[13] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[14] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[15] ), 
            .O(n7479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11380.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11381 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[11] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[18] ), 
            .I2(n7479), .O(n7480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11381.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11382 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[20] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[21] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[22] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[23] ), 
            .O(n7481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11382.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11383 (.I0(n7478), .I1(n7480), .I2(n7481), .O(n7482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11383.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11384 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[0] ), 
            .I1(n1642), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11384.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11385 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[21] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[22] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[23] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[24] ), 
            .O(n7483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11385.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11386 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[17] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[18] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[19] ), 
            .I3(n7483), .O(n7484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11386.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11387 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[13] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[14] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[15] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[16] ), 
            .O(n7485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11387.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11388 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[20] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[25] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[26] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[27] ), 
            .O(n7486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11388.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11389 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[11] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[12] ), 
            .I2(n7485), .I3(n7486), .O(n7487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11389.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11390 (.I0(n7484), .I1(n7487), .O(n7488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11390.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11391 (.I0(DdrCtrl_ALEN_0[0]), .I1(n1473), .I2(n7488), 
            .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11391.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11392 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcx_location[10] ), 
            .I1(n1471), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11392.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11393 (.I0(n1640), .I1(n1469), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n333 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11393.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11394 (.I0(n1359), .I1(n1467), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11394.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11395 (.I0(n1357), .I1(n1465), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11395.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11396 (.I0(n1355), .I1(n1463), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11396.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11397 (.I0(n1353), .I1(n1461), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n329 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11397.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11398 (.I0(n1351), .I1(n1459), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11398.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11399 (.I0(n1327), .I1(n1457), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n327 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11399.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11400 (.I0(n1325), .I1(n1455), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11400.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11401 (.I0(n1323), .I1(n1453), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11401.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11402 (.I0(n1321), .I1(n1451), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11402.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11403 (.I0(n1319), .I1(n1449), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n323 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11403.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11404 (.I0(n1317), .I1(n1405), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11404.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11405 (.I0(n1315), .I1(n1403), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n321 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11405.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11406 (.I0(n1313), .I1(n1401), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11406.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11407 (.I0(n1311), .I1(n1399), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11407.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11408 (.I0(n1309), .I1(n1397), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11408.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11409 (.I0(n1308), .I1(n1396), .I2(n7488), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11409.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11410 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[1] ), 
            .I1(n1306), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11410.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11411 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[2] ), 
            .I1(n1304), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11411.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11412 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[3] ), 
            .I1(n1302), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11412.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11413 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[4] ), 
            .I1(n1300), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11413.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11414 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[5] ), 
            .I1(n1298), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11414.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11415 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[6] ), 
            .I1(n1296), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11415.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11416 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[7] ), 
            .I1(n1294), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11416.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11417 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[8] ), 
            .I1(n1292), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11417.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11418 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[9] ), 
            .I1(n1290), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11418.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11419 (.I0(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/genblk1.temp_srcy_location[10] ), 
            .I1(n1288), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11419.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11420 (.I0(n1672), .I1(n1286), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11420.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11421 (.I0(n1249), .I1(n1284), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11421.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11422 (.I0(n1247), .I1(n1282), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11422.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11423 (.I0(n1245), .I1(n1280), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11423.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11424 (.I0(n1243), .I1(n1278), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11424.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11425 (.I0(n1241), .I1(n1276), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11425.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11426 (.I0(n1239), .I1(n1274), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11426.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11427 (.I0(n1237), .I1(n1272), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11427.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11428 (.I0(n1235), .I1(n1266), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11428.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11429 (.I0(n1233), .I1(n1264), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11429.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11430 (.I0(n1231), .I1(n1262), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11430.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11431 (.I0(n1229), .I1(n1260), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11431.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11432 (.I0(n1227), .I1(n1258), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11432.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11433 (.I0(n1225), .I1(n1256), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11433.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11434 (.I0(n1223), .I1(n1254), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11434.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11435 (.I0(n1221), .I1(n1252), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11435.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11436 (.I0(n1220), .I1(n1251), .I2(n7482), .O(\u_scaler_gray/u1_bilinear_gray/u0_cal_bilinear_srcxy/n435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11436.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11437 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21] ), 
            .O(n7489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11437.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11438 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15] ), 
            .I2(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17] ), 
            .O(n7490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11438.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11439 (.I0(n7489), .I1(n7490), .I2(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12] ), 
            .I3(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13] ), 
            .O(n7491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11439.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11440 (.I0(n7491), .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[11] ), 
            .O(n7492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11440.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11441 (.I0(n7492), .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[12] ), 
            .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11441.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11442 (.I0(DdrCtrl_WVALID_0), .I1(DdrCtrl_WREADY_0), .O(\u_axi4_ctrl/n363 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11442.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11443 (.I0(n653), .I1(n655), .I2(n657), .I3(n2355), 
            .O(n7493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11443.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11444 (.I0(n645), .I1(n647), .I2(n649), .I3(n651), 
            .O(n7494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11444.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11445 (.I0(n642), .I1(n643), .I2(n7493), .I3(n7494), 
            .O(n7495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11445.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11446 (.I0(\u_axi4_ctrl/wfifo_empty ), .I1(\u_axi4_ctrl/n363 ), 
            .I2(n7495), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__11446.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__11447 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), .O(n7496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11447.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11448 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] ), 
            .O(n7497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11448.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11449 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
            .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .O(n7498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0990 */ ;
    defparam LUT__11449.LUTMASK = 16'h0990;
    EFX_LUT4 LUT__11450 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .I2(n7497), .I3(n7498), .O(n7499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__11450.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__11451 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .O(n7500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11451.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11452 (.I0(n7499), .I1(n7500), .I2(n7496), .I3(tvalid_o), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__11452.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__11453 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[8] ), 
            .I1(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/round_data[9] ), 
            .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n357 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__11453.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__11454 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[13] ), 
            .I1(n1913), .I2(n7492), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n343 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11454.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11455 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[14] ), 
            .I1(n936), .I2(n7492), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11455.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11456 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[15] ), 
            .I1(n932), .I2(n7492), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n341 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11456.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11457 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[16] ), 
            .I1(n930), .I2(n7492), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11457.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11458 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[17] ), 
            .I1(n926), .I2(n7492), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n339 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11458.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11459 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[18] ), 
            .I1(n924), .I2(n7492), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11459.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11460 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[19] ), 
            .I1(n922), .I2(n7492), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n337 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11460.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11461 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[20] ), 
            .I1(n920), .I2(n7492), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11461.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11462 (.I0(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/level2_add0[21] ), 
            .I1(n919), .I2(n7492), .O(\u_scaler_gray/u1_bilinear_gray/u2_cal_bilinear_data/n335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11462.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11463 (.I0(\u_axi4_ctrl/wframe_index[1] ), .I1(\u_axi4_ctrl/wframe_index[0] ), 
            .O(\u_axi4_ctrl/n316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11463.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11464 (.I0(\u_axi4_ctrl/wframe_vsync_dly[2] ), .I1(\u_axi4_ctrl/wframe_vsync_dly[3] ), 
            .O(\u_axi4_ctrl/equal_38/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11464.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11468 (.I0(\u_axi4_ctrl/wframe_vsync_dly[3] ), .I1(\u_axi4_ctrl/wframe_vsync_dly[2] ), 
            .I2(\Axi0ResetReg[2] ), .O(\u_axi4_ctrl/n1469 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__11468.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__11469 (.I0(\u_axi4_ctrl/wframe_index[1] ), .I1(\u_axi4_ctrl/wframe_index[0] ), 
            .O(\u_axi4_ctrl/n317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11469.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11470 (.I0(\u_axi4_ctrl/wframe_index[0] ), .I1(\u_axi4_ctrl/wframe_index[1] ), 
            .O(\u_axi4_ctrl/n336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11470.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11471 (.I0(\u_axi4_ctrl/rframe_vsync_dly[2] ), .I1(\u_axi4_ctrl/rframe_vsync_dly[3] ), 
            .O(\u_axi4_ctrl/equal_47/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11471.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11472 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/rdata_cnt_dly[3] ), 
            .O(n7503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11472.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11473 (.I0(n7503), .I1(\u_axi4_ctrl/rdata_cnt_dly[4] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[5] ), .O(n7504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11473.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11474 (.I0(DdrCtrl_RREADY_0), .I1(DdrCtrl_RVALID_0), .O(\u_axi4_ctrl/n379 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11474.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11475 (.I0(\u_axi4_ctrl/rdata_cnt_dly[7] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[8] ), 
            .I2(\u_axi4_ctrl/n379 ), .O(n7505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11475.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11476 (.I0(\u_axi4_ctrl/rdata_cnt_dly[6] ), .I1(n7504), 
            .I2(n7505), .O(\u_axi4_ctrl/n381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11476.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11477 (.I0(\u_axi4_ctrl/n381 ), .I1(\u_axi4_ctrl/state[1] ), 
            .I2(\u_axi4_ctrl/state[2] ), .O(n7506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__11477.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__11478 (.I0(DdrCtrl_BVALID_0), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(DdrCtrl_WREADY_0), .I3(n7041), .O(n7507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__11478.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__11479 (.I0(n426), .I1(n428), .I2(n430), .I3(n2520), 
            .O(n7508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11479.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11480 (.I0(n422), .I1(n424), .I2(n7508), .I3(n420), 
            .O(n7509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__11480.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__11481 (.I0(n7509), .I1(n419), .O(n7510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11481.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11482 (.I0(n557), .I1(n558), .O(n7511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11482.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11483 (.I0(n7511), .I1(n7510), .I2(DdrCtrl_AREADY_0), 
            .I3(\u_axi4_ctrl/state[0] ), .O(n7512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__11483.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__11484 (.I0(n7512), .I1(n7507), .I2(\u_axi4_ctrl/state[2] ), 
            .I3(\u_axi4_ctrl/state[1] ), .O(n7513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__11484.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__11485 (.I0(DdrCtrl_AREADY_0), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(n7506), .I3(n7513), .O(\u_axi4_ctrl/n389 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0 */ ;
    defparam LUT__11485.LUTMASK = 16'hffe0;
    EFX_LUT4 LUT__11486 (.I0(n7511), .I1(\u_axi4_ctrl/state[0] ), .I2(\u_axi4_ctrl/state[1] ), 
            .I3(\u_axi4_ctrl/state[2] ), .O(\u_axi4_ctrl/n405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11486.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11487 (.I0(\u_axi4_ctrl/state[0] ), .I1(\u_axi4_ctrl/state[1] ), 
            .I2(\u_axi4_ctrl/state[2] ), .I3(n7510), .O(n7514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11487.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11488 (.I0(n7514), .I1(\Axi0ResetReg[2] ), .O(\u_axi4_ctrl/n1476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11488.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11489 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .O(n7515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11489.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11490 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .O(n7516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11490.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11491 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] ), 
            .I2(n7515), .I3(n7516), .O(n7517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__11491.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__11492 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), .O(n7518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11492.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11493 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .O(n7519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11493.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11494 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .O(n7520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11494.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11495 (.I0(n7518), .I1(n7519), .I2(n7517), .I3(n7520), 
            .O(n7521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11495.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11496 (.I0(lcd_de), .I1(\u_axi4_ctrl/rfifo_empty ), .I2(n7521), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__11496.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__11497 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] ), 
            .O(n7522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11497.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11498 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .O(n7523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11498.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11499 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[12] ), 
            .O(n7524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0990 */ ;
    defparam LUT__11499.LUTMASK = 16'h0990;
    EFX_LUT4 LUT__11500 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] ), 
            .I2(n7523), .I3(n7524), .O(n7525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__11500.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__11501 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] ), 
            .O(n7526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__11501.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__11502 (.I0(n7525), .I1(n7526), .I2(n7522), .I3(\u_axi4_ctrl/rfifo_wenb ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__11502.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__11505 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .O(\u_axi4_ctrl/n1544 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11505.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11508 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
            .I1(\u_axi4_ctrl/n363 ), .O(ceg_net289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11508.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11509 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11509.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11510 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11510.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11511 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11511.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11512 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11512.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11513 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11513.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11514 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11514.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11515 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11515.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11516 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11516.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11517 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), .I2(\u_axi4_ctrl/wfifo_empty ), 
            .O(n5870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11517.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11518 (.I0(n4225), .I1(n5870), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11518.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11521 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11521.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11522 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11522.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11523 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11523.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11524 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11524.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11525 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11525.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11526 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11526.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11527 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11527.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11528 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11528.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11529 (.I0(n4222), .I1(n4225), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11529.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11530 (.I0(n4211), .I1(n4222), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11530.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11531 (.I0(n4176), .I1(n4211), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11531.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11532 (.I0(n4138), .I1(n4176), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11532.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11533 (.I0(n4135), .I1(n4138), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11533.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11534 (.I0(n4132), .I1(n4135), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11534.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11535 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[8] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11535.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11536 (.I0(n4132), .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[8] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11536.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11537 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11537.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11538 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11538.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11539 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11539.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11540 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11540.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11541 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11541.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11542 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11542.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11543 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11543.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11544 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11544.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11545 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
            .I1(lcd_de), .O(ceg_net296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11545.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11546 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11546.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11547 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11547.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11548 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11548.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11549 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11549.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11550 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11550.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11551 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11551.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11552 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11552.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11553 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11553.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11554 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11554.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11557 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[12] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11557.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11558 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[11] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11558.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11559 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11559.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11560 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11560.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11561 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11561.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11562 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11562.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11563 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11563.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11564 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11564.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11565 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .O(n7527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11565.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11566 (.I0(n7527), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11566.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11567 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .O(n7528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11567.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11568 (.I0(n7528), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11568.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11569 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .O(n7529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11569.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11570 (.I0(n7529), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11570.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11571 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .O(n7530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11571.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11572 (.I0(n7530), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11572.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11573 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .O(n7531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11573.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11574 (.I0(n7531), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11574.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11575 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] ), 
            .O(n7532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11575.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11576 (.I0(n7532), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11576.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11577 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[11] ), .I2(\u_axi4_ctrl/rfifo_empty ), 
            .O(n7533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11577.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11578 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] ), 
            .I2(\u_axi4_ctrl/rfifo_empty ), .I3(n7533), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53 */ ;
    defparam LUT__11578.LUTMASK = 16'hac53;
    EFX_LUT4 LUT__11579 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[12] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[12] ), 
            .I2(\u_axi4_ctrl/rfifo_empty ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11579.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11580 (.I0(n7533), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[12] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11580.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11581 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11581.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11582 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11582.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11583 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11583.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11584 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11584.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11585 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11585.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11586 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11586.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11587 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11587.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11588 (.I0(\u_axi4_ctrl/wframe_index[1] ), .I1(\u_axi4_ctrl/wframe_index[0] ), 
            .O(\u_axi4_ctrl/n335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11588.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11589 (.I0(\u_axi4_ctrl/state[2] ), .I1(\u_axi4_ctrl/state[0] ), 
            .O(n7534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11589.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11590 (.I0(DdrCtrl_AREADY_0), .I1(DdrCtrl_BVALID_0), .I2(n7534), 
            .I3(\u_axi4_ctrl/state[1] ), .O(\u_axi4_ctrl/n1610 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3fa0 */ ;
    defparam LUT__11590.LUTMASK = 16'h3fa0;
    EFX_LUT4 LUT__11591 (.I0(\u_axi4_ctrl/state[2] ), .I1(\Axi0ResetReg[2] ), 
            .O(\u_axi4_ctrl/n1617 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__11591.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__11592 (.I0(n7506), .I1(n7514), .O(\u_axi4_ctrl/n387 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__11592.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__11593 (.I0(DdrCtrl_BREADY_0), .I1(DdrCtrl_BVALID_0), .O(\u_axi4_ctrl/n369 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11593.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11594 (.I0(n6320), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .O(n6323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11594.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11595 (.I0(n6326), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .O(n6329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11595.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11596 (.I0(n6332), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .O(n6335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11596.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11597 (.I0(n6335), .I1(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] ), 
            .O(n6338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11597.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11598 (.I0(\u_axi4_ctrl/rframe_vsync_dly[3] ), .I1(\u_axi4_ctrl/rframe_vsync_dly[2] ), 
            .I2(\Axi0ResetReg[2] ), .O(\u_axi4_ctrl/n1478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__11598.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__11599 (.I0(\u_axi4_ctrl/awaddr[10] ), .I1(\u_axi4_ctrl/araddr[10] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11599.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11600 (.I0(\u_axi4_ctrl/n1476 ), .I1(\u_axi4_ctrl/n405 ), 
            .O(ceg_net401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11600.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11601 (.I0(\u_axi4_ctrl/awaddr[11] ), .I1(\u_axi4_ctrl/araddr[11] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11601.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11602 (.I0(\u_axi4_ctrl/awaddr[12] ), .I1(\u_axi4_ctrl/araddr[12] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n695 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11602.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11603 (.I0(\u_axi4_ctrl/awaddr[13] ), .I1(\u_axi4_ctrl/araddr[13] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11603.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11604 (.I0(\u_axi4_ctrl/awaddr[14] ), .I1(\u_axi4_ctrl/araddr[14] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11604.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11605 (.I0(\u_axi4_ctrl/awaddr[15] ), .I1(\u_axi4_ctrl/araddr[15] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11605.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11606 (.I0(\u_axi4_ctrl/awaddr[16] ), .I1(\u_axi4_ctrl/araddr[16] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11606.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11607 (.I0(\u_axi4_ctrl/awaddr[17] ), .I1(\u_axi4_ctrl/araddr[17] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11607.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11608 (.I0(\u_axi4_ctrl/awaddr[18] ), .I1(\u_axi4_ctrl/araddr[18] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n689 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11608.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11609 (.I0(\u_axi4_ctrl/awaddr[19] ), .I1(\u_axi4_ctrl/araddr[19] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n688 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11609.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11610 (.I0(\u_axi4_ctrl/awaddr[20] ), .I1(\u_axi4_ctrl/araddr[20] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n687 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11610.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11611 (.I0(\u_axi4_ctrl/awaddr[21] ), .I1(\u_axi4_ctrl/araddr[21] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n686 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11611.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11612 (.I0(\u_axi4_ctrl/awaddr[22] ), .I1(\u_axi4_ctrl/araddr[22] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n685 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11612.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11613 (.I0(\u_axi4_ctrl/awaddr[23] ), .I1(\u_axi4_ctrl/araddr[23] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11613.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11614 (.I0(\u_axi4_ctrl/wframe_index[0] ), .I1(\u_axi4_ctrl/rframe_index[0] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n683 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11614.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11615 (.I0(\u_axi4_ctrl/wframe_index[1] ), .I1(\u_axi4_ctrl/rframe_index[1] ), 
            .I2(n7514), .O(\u_axi4_ctrl/n682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11615.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11616 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .O(\u_axi4_ctrl/n1499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11616.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11617 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .O(\u_axi4_ctrl/n1504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11617.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11618 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/wdata_cnt_dly[3] ), 
            .O(\u_axi4_ctrl/n1509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11618.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11619 (.I0(n7038), .I1(\u_axi4_ctrl/wdata_cnt_dly[4] ), 
            .O(\u_axi4_ctrl/n1514 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11619.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11620 (.I0(n7038), .I1(\u_axi4_ctrl/wdata_cnt_dly[4] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[5] ), .O(\u_axi4_ctrl/n1519 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11620.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11621 (.I0(n7039), .I1(\u_axi4_ctrl/wdata_cnt_dly[6] ), 
            .O(\u_axi4_ctrl/n1524 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11621.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11622 (.I0(n7039), .I1(\u_axi4_ctrl/wdata_cnt_dly[6] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[7] ), .O(\u_axi4_ctrl/n1529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11622.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11623 (.I0(n7039), .I1(\u_axi4_ctrl/wdata_cnt_dly[6] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[7] ), .I3(\u_axi4_ctrl/wdata_cnt_dly[8] ), 
            .O(\u_axi4_ctrl/n1534 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11623.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11624 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[2] ), .O(\u_axi4_ctrl/n1549 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11624.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11625 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/rdata_cnt_dly[3] ), 
            .O(\u_axi4_ctrl/n1554 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11625.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11626 (.I0(n7503), .I1(\u_axi4_ctrl/rdata_cnt_dly[4] ), 
            .O(\u_axi4_ctrl/n1559 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11626.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11627 (.I0(n7503), .I1(\u_axi4_ctrl/rdata_cnt_dly[4] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[5] ), .O(\u_axi4_ctrl/n1564 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11627.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11628 (.I0(n7504), .I1(\u_axi4_ctrl/rdata_cnt_dly[6] ), 
            .O(\u_axi4_ctrl/n1569 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__11628.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__11629 (.I0(n7504), .I1(\u_axi4_ctrl/rdata_cnt_dly[6] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[7] ), .O(\u_axi4_ctrl/n1574 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11629.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11630 (.I0(n7504), .I1(\u_axi4_ctrl/rdata_cnt_dly[6] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[7] ), .I3(\u_axi4_ctrl/rdata_cnt_dly[8] ), 
            .O(\u_axi4_ctrl/n1579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__11630.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__11631 (.I0(\u_lcd_driver/vcnt[1] ), .I1(\u_lcd_driver/vcnt[2] ), 
            .O(n7535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11631.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11632 (.I0(\u_lcd_driver/vcnt[3] ), .I1(\u_lcd_driver/vcnt[4] ), 
            .I2(\u_lcd_driver/vcnt[5] ), .I3(\u_lcd_driver/vcnt[6] ), .O(n7536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11632.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11633 (.I0(n7536), .I1(n7535), .I2(\u_lcd_driver/vcnt[7] ), 
            .I3(\u_lcd_driver/vcnt[8] ), .O(n7537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__11633.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__11634 (.I0(\u_lcd_driver/vcnt[9] ), .I1(n7537), .I2(\u_lcd_driver/vcnt[10] ), 
            .I3(\u_lcd_driver/vcnt[11] ), .O(n7538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__11634.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__11635 (.I0(\u_lcd_driver/vcnt[0] ), .I1(n7538), .O(\u_lcd_driver/n83 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11635.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11636 (.I0(\u_lcd_driver/hcnt[0] ), .I1(\u_lcd_driver/hcnt[1] ), 
            .I2(\u_lcd_driver/hcnt[2] ), .I3(\u_lcd_driver/hcnt[3] ), .O(n7539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__11636.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__11637 (.I0(n7539), .I1(\u_lcd_driver/hcnt[4] ), .I2(\u_lcd_driver/hcnt[5] ), 
            .O(n7540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11637.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11638 (.I0(\u_lcd_driver/hcnt[6] ), .I1(\u_lcd_driver/hcnt[7] ), 
            .I2(\u_lcd_driver/hcnt[9] ), .I3(\u_lcd_driver/hcnt[11] ), .O(n7541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11638.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11639 (.I0(n7540), .I1(n7541), .I2(\u_lcd_driver/hcnt[8] ), 
            .I3(\u_lcd_driver/hcnt[10] ), .O(\u_lcd_driver/equal_17/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__11639.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__11640 (.I0(\u_lcd_driver/hcnt[4] ), .I1(\u_lcd_driver/hcnt[3] ), 
            .I2(\u_lcd_driver/hcnt[5] ), .I3(\u_lcd_driver/hcnt[8] ), .O(n7542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__11640.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__11641 (.I0(\u_lcd_driver/hcnt[10] ), .I1(n7542), .I2(n7541), 
            .O(\u_lcd_driver/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__11641.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__11642 (.I0(\u_lcd_driver/vcnt[2] ), .I1(\u_lcd_driver/vcnt[3] ), 
            .I2(\u_lcd_driver/vcnt[4] ), .I3(\u_lcd_driver/vcnt[5] ), .O(n7543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11642.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11643 (.I0(\u_lcd_driver/vcnt[1] ), .I1(\u_lcd_driver/vcnt[0] ), 
            .I2(n7543), .O(n7544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__11643.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__11644 (.I0(\u_lcd_driver/vcnt[6] ), .I1(\u_lcd_driver/vcnt[7] ), 
            .I2(\u_lcd_driver/vcnt[8] ), .I3(\u_lcd_driver/vcnt[9] ), .O(n7545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__11644.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__11645 (.I0(\u_lcd_driver/vcnt[10] ), .I1(\u_lcd_driver/vcnt[11] ), 
            .I2(n7544), .I3(n7545), .O(\u_lcd_driver/n97 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__11645.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__11646 (.I0(\u_lcd_driver/vcnt[0] ), .I1(\u_lcd_driver/vcnt[1] ), 
            .I2(\u_lcd_driver/vcnt[2] ), .O(n7546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__11646.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__11647 (.I0(n7546), .I1(\u_lcd_driver/vcnt[3] ), .I2(\u_lcd_driver/vcnt[4] ), 
            .I3(\u_lcd_driver/vcnt[5] ), .O(n7547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h07e0 */ ;
    defparam LUT__11647.LUTMASK = 16'h07e0;
    EFX_LUT4 LUT__11648 (.I0(n7545), .I1(\u_lcd_driver/vcnt[6] ), .I2(n7547), 
            .I3(\u_lcd_driver/vcnt[5] ), .O(n7548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__11648.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__11649 (.I0(\u_lcd_driver/vcnt[7] ), .I1(\u_lcd_driver/vcnt[8] ), 
            .I2(n7548), .I3(\u_lcd_driver/vcnt[9] ), .O(n7549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__11649.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__11650 (.I0(\u_lcd_driver/hcnt[6] ), .I1(\u_lcd_driver/hcnt[5] ), 
            .I2(\u_lcd_driver/hcnt[7] ), .O(n7550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__11650.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__11651 (.I0(n7550), .I1(\u_lcd_driver/hcnt[8] ), .I2(\u_lcd_driver/hcnt[9] ), 
            .I3(\u_lcd_driver/hcnt[10] ), .O(n7551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h01fe */ ;
    defparam LUT__11651.LUTMASK = 16'h01fe;
    EFX_LUT4 LUT__11652 (.I0(\u_lcd_driver/vcnt[10] ), .I1(\u_lcd_driver/vcnt[11] ), 
            .I2(\u_lcd_driver/hcnt[11] ), .I3(n7551), .O(n7552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__11652.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__11653 (.I0(\u_lcd_driver/vcnt[5] ), .I1(n7548), .I2(n7549), 
            .I3(n7552), .O(\u_lcd_driver/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__11653.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__11654 (.I0(\u_lcd_driver/vcnt[6] ), .I1(n7544), .I2(\u_lcd_driver/vcnt[7] ), 
            .I3(\u_lcd_driver/vcnt[8] ), .O(n7553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__11654.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__11655 (.I0(n7553), .I1(\u_lcd_driver/vcnt[9] ), .I2(n7552), 
            .O(\u_lcd_driver/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__11655.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__11656 (.I0(\u_lcd_driver/hcnt[9] ), .I1(\u_lcd_driver/hcnt[8] ), 
            .I2(\u_lcd_driver/hcnt[10] ), .I3(\u_lcd_driver/hcnt[11] ), 
            .O(n7554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__11656.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__11657 (.I0(n7541), .I1(n7540), .I2(n7554), .O(n7555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__11657.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__11658 (.I0(n7555), .I1(\u_lcd_driver/hcnt[0] ), .O(\u_lcd_driver/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__11658.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__11659 (.I0(n7538), .I1(n3029), .O(\u_lcd_driver/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11659.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11660 (.I0(n7538), .I1(n398), .O(\u_lcd_driver/n81 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11660.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11661 (.I0(n7538), .I1(n396), .O(\u_lcd_driver/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11661.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11662 (.I0(n7538), .I1(n394), .O(\u_lcd_driver/n79 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11662.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11663 (.I0(n7538), .I1(n392), .O(\u_lcd_driver/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11663.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11664 (.I0(n7538), .I1(n390), .O(\u_lcd_driver/n77 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11664.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11665 (.I0(n7538), .I1(n388), .O(\u_lcd_driver/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11665.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11666 (.I0(n7538), .I1(n386), .O(\u_lcd_driver/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11666.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11667 (.I0(n7538), .I1(n384), .O(\u_lcd_driver/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11667.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11668 (.I0(n7538), .I1(n382), .O(\u_lcd_driver/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11668.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11669 (.I0(n7538), .I1(n381), .O(\u_lcd_driver/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__11669.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__11670 (.I0(n7555), .I1(n2537), .O(\u_lcd_driver/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11670.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11671 (.I0(n7555), .I1(n417), .O(\u_lcd_driver/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11671.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11672 (.I0(n7555), .I1(n415), .O(\u_lcd_driver/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11672.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11673 (.I0(n7555), .I1(n413), .O(\u_lcd_driver/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11673.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11674 (.I0(n7555), .I1(n411), .O(\u_lcd_driver/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11674.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11675 (.I0(n7555), .I1(n409), .O(\u_lcd_driver/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11675.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11676 (.I0(n7555), .I1(n407), .O(\u_lcd_driver/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11676.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11677 (.I0(n7555), .I1(n405), .O(\u_lcd_driver/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11677.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11678 (.I0(n7555), .I1(n403), .O(\u_lcd_driver/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11678.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11679 (.I0(n7555), .I1(n401), .O(\u_lcd_driver/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11679.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11680 (.I0(n7555), .I1(n400), .O(\u_lcd_driver/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__11680.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__11681 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I1(n7375), .I2(n7378), .I3(n7353), .O(n7556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc531 */ ;
    defparam LUT__11681.LUTMASK = 16'hc531;
    EFX_LUT4 LUT__11682 (.I0(lcd_hs), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q ), 
            .I2(n7556), .I3(lcd_de), .O(\u_rgb2dvi/enc_0/n869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3aa */ ;
    defparam LUT__11682.LUTMASK = 16'hc3aa;
    EFX_LUT4 LUT__11683 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_19_q ), .O(n7557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11683.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11684 (.I0(lcd_hs), .I1(n7557), .I2(n7556), .I3(lcd_de), 
            .O(\u_rgb2dvi/enc_0/n764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11684.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11685 (.I0(lcd_hs), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21_q ), 
            .I2(n7556), .I3(lcd_de), .O(\u_rgb2dvi/enc_0/n770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__11685.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__11686 (.I0(lcd_hs), .I1(n7556), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18_q ), 
            .I3(lcd_de), .O(\u_rgb2dvi/enc_0/n776 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3aa */ ;
    defparam LUT__11686.LUTMASK = 16'hc3aa;
    EFX_LUT4 LUT__11687 (.I0(lcd_hs), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_q ), 
            .I2(n7556), .I3(lcd_de), .O(\u_rgb2dvi/enc_0/n782 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__11687.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__11688 (.I0(\u_lcd_driver/r_lcd_dv ), .I1(\u_lcd_driver/r_lcd_rgb[5] ), 
            .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_q ), .O(n7558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__11688.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__11689 (.I0(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I1(n7558), .O(n7559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__11689.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__11690 (.I0(lcd_hs), .I1(n7559), .I2(n7556), .I3(lcd_de), 
            .O(\u_rgb2dvi/enc_0/n788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11690.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11691 (.I0(lcd_hs), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25_q ), 
            .I2(n7556), .I3(lcd_de), .O(\u_rgb2dvi/enc_0/n794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc355 */ ;
    defparam LUT__11691.LUTMASK = 16'hc355;
    EFX_LUT4 LUT__11692 (.I0(lcd_hs), .I1(n7341), .I2(n7556), .I3(lcd_de), 
            .O(\u_rgb2dvi/enc_0/n800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3caa */ ;
    defparam LUT__11692.LUTMASK = 16'h3caa;
    EFX_LUT4 LUT__11693 (.I0(lcd_hs), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(lcd_de), .O(\u_rgb2dvi/enc_0/n806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__11693.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__11694 (.I0(n7556), .I1(lcd_hs), .I2(lcd_vs), .I3(lcd_de), 
            .O(\u_rgb2dvi/enc_0/n812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h55c3 */ ;
    defparam LUT__11694.LUTMASK = 16'h55c3;
    EFX_LUT4 LUT__11695 (.I0(n7368), .I1(n7366), .I2(n7353), .O(n7560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__11695.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__11696 (.I0(n7368), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7560), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q ), .O(\u_rgb2dvi/enc_1/q_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f */ ;
    defparam LUT__11696.LUTMASK = 16'hb04f;
    EFX_LUT4 LUT__11697 (.I0(n7368), .I1(n7560), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_19_q ), 
            .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .O(\u_rgb2dvi/enc_1/q_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h78c3 */ ;
    defparam LUT__11697.LUTMASK = 16'h78c3;
    EFX_LUT4 LUT__11698 (.I0(n7368), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7560), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21_q ), 
            .O(\u_rgb2dvi/enc_1/q_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f */ ;
    defparam LUT__11698.LUTMASK = 16'hb04f;
    EFX_LUT4 LUT__11699 (.I0(n7368), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7560), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18_q ), 
            .O(\u_rgb2dvi/enc_1/q_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f */ ;
    defparam LUT__11699.LUTMASK = 16'hb04f;
    EFX_LUT4 LUT__11700 (.I0(n7368), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7560), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_q ), 
            .O(\u_rgb2dvi/enc_1/q_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f */ ;
    defparam LUT__11700.LUTMASK = 16'hb04f;
    EFX_LUT4 LUT__11701 (.I0(n7368), .I1(n7560), .I2(n7558), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .O(\u_rgb2dvi/enc_1/q_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h78c3 */ ;
    defparam LUT__11701.LUTMASK = 16'h78c3;
    EFX_LUT4 LUT__11702 (.I0(n7368), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7560), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25_q ), 
            .O(\u_rgb2dvi/enc_1/q_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f */ ;
    defparam LUT__11702.LUTMASK = 16'hb04f;
    EFX_LUT4 LUT__11703 (.I0(n7368), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7560), .I3(n7341), .O(\u_rgb2dvi/enc_1/q_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4fb0 */ ;
    defparam LUT__11703.LUTMASK = 16'h4fb0;
    EFX_LUT4 LUT__11704 (.I0(n7368), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7560), .O(\u_rgb2dvi/enc_1/q_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__11704.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__11705 (.I0(n7358), .I1(n7325), .I2(n7353), .O(n7561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__11705.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__11706 (.I0(n7358), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7561), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q ), .O(\u_rgb2dvi/enc_2/q_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f */ ;
    defparam LUT__11706.LUTMASK = 16'hb04f;
    EFX_LUT4 LUT__11707 (.I0(n7358), .I1(n7561), .I2(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_19_q ), 
            .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .O(\u_rgb2dvi/enc_2/q_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h78c3 */ ;
    defparam LUT__11707.LUTMASK = 16'h78c3;
    EFX_LUT4 LUT__11708 (.I0(n7358), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7561), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21_q ), 
            .O(\u_rgb2dvi/enc_2/q_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f */ ;
    defparam LUT__11708.LUTMASK = 16'hb04f;
    EFX_LUT4 LUT__11709 (.I0(n7358), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7561), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18_q ), 
            .O(\u_rgb2dvi/enc_2/q_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f */ ;
    defparam LUT__11709.LUTMASK = 16'hb04f;
    EFX_LUT4 LUT__11710 (.I0(n7358), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7561), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_q ), 
            .O(\u_rgb2dvi/enc_2/q_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f */ ;
    defparam LUT__11710.LUTMASK = 16'hb04f;
    EFX_LUT4 LUT__11711 (.I0(n7358), .I1(n7561), .I2(n7558), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .O(\u_rgb2dvi/enc_2/q_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h78c3 */ ;
    defparam LUT__11711.LUTMASK = 16'h78c3;
    EFX_LUT4 LUT__11712 (.I0(n7358), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7561), .I3(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25_q ), 
            .O(\u_rgb2dvi/enc_2/q_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb04f */ ;
    defparam LUT__11712.LUTMASK = 16'hb04f;
    EFX_LUT4 LUT__11713 (.I0(n7358), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7561), .I3(n7341), .O(\u_rgb2dvi/enc_2/q_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4fb0 */ ;
    defparam LUT__11713.LUTMASK = 16'h4fb0;
    EFX_LUT4 LUT__11714 (.I0(n7358), .I1(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q ), 
            .I2(n7561), .O(\u_rgb2dvi/enc_2/q_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__11714.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__11715 (.I0(\r_hdmi_tx0_o[6] ), .I1(\w_hdmi_txd0[1] ), 
            .I2(rc_hdmi_tx), .O(n591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11715.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11716 (.I0(\r_hdmi_tx0_o[7] ), .I1(\w_hdmi_txd0[2] ), 
            .I2(rc_hdmi_tx), .O(n590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__11716.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__11717 (.I0(\r_hdmi_tx0_o[8] ), .I1(\w_hdmi_txd0[3] ), 
            .I2(rc_hdmi_tx), .O(n589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11717.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11718 (.I0(\r_hdmi_tx0_o[9] ), .I1(\w_hdmi_txd0[4] ), 
            .I2(rc_hdmi_tx), .O(n588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__11718.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__11719 (.I0(\r_hdmi_tx1_o[6] ), .I1(\w_hdmi_txd1[1] ), 
            .I2(rc_hdmi_tx), .O(n602_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11719.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11720 (.I0(\r_hdmi_tx1_o[7] ), .I1(\w_hdmi_txd1[2] ), 
            .I2(rc_hdmi_tx), .O(n601_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__11720.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__11721 (.I0(\r_hdmi_tx1_o[8] ), .I1(\w_hdmi_txd1[3] ), 
            .I2(rc_hdmi_tx), .O(n600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11721.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11722 (.I0(\r_hdmi_tx1_o[9] ), .I1(\w_hdmi_txd1[4] ), 
            .I2(rc_hdmi_tx), .O(n599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__11722.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__11723 (.I0(\r_hdmi_tx2_o[6] ), .I1(\w_hdmi_txd2[1] ), 
            .I2(rc_hdmi_tx), .O(n613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11723.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11724 (.I0(\r_hdmi_tx2_o[7] ), .I1(\w_hdmi_txd2[2] ), 
            .I2(rc_hdmi_tx), .O(n612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__11724.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__11725 (.I0(\r_hdmi_tx1_o[8] ), .I1(\w_hdmi_txd2[3] ), 
            .I2(rc_hdmi_tx), .O(n611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__11725.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__11726 (.I0(\r_hdmi_tx2_o[9] ), .I1(\w_hdmi_txd2[4] ), 
            .I2(rc_hdmi_tx), .O(n610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__11726.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__11811 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
            .O(DdrCtrl_CFG_SEQ_RST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11811.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11835 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[0] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[0]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11835.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11836 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[1] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[1]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11836.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11837 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[2] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[2]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11837.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11838 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[3] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[3]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11838.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11839 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[4] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[4]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11839.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11840 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[5] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[5]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11840.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11841 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[6] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[6]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11841.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11842 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[7] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[7]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11842.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11843 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[8] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[8]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11843.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11844 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[9] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[9]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11844.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11845 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[10]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11845.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11846 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb00[11]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11846.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11848 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[0] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[0]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11848.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11849 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[1] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[1]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11849.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11850 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[2] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[2]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11850.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11851 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[3] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[3]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11851.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11852 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[4] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[4]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11852.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11853 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[5] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[5]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11853.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11854 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[6] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[6]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11854.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11855 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[7] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[7]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11855.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11856 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[8] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[8]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11856.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11857 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[9] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[9]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11857.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11858 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[10]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11858.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11859 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb01[11]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11859.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11860 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[8] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[8]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11860.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11861 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[9] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[9]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11861.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11862 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[10]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11862.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11863 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb10[11]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11863.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11864 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[8] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[8]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11864.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11865 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[9] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[9]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11865.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11866 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[10] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[10]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11866.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__11867 (.I0(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11] ), 
            .O(\u_scaler_gray/u0_data_stream_ctr/r_addrb11[11]__I )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__11867.LUTMASK = 16'h5555;
    EFX_FF \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26  (.D(n6895), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[1]~FF_frt_13_frt_26 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25  (.D(n7340), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_25 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24  (.D(n7349), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_24 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[5]~FF_frt_23  (.D(n7350), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[5]~FF_frt_23_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_23 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_23 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_23 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_23 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_23 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_23 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[5]~FF_frt_23 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12  (.D(n7328), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21  (.D(n7343), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_21 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_19  (.D(n7344), .CE(1'b1), 
           .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_19_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_19 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_19 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_19 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_19 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_19 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_19 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_19 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18  (.D(n7347), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_12_frt_17_frt_18 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20  (.D(\u_rgb2dvi/enc_0/n103 ), 
           .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_3_frt_11_frt_16_frt_20 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_dv~FF_frt_7  (.D(n7335), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\u_lcd_driver/r_lcd_dv~FF_frt_7_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_dv~FF_frt_7 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4  (.D(n7333), .CE(1'b1), .CLK(\hdmi_clk1x_i~O ), 
           .SR(1'b0), .Q(\u_lcd_driver/r_lcd_rgb[0]~FF_frt_4_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, INIT_VALUE=1'b0 */ ;   // C:\Users\Yuanbing Ouyang\Desktop\xidianFPGA\T35\scale\01efx_bilinear_scaler_hdmi\ar0135_dvp_lvds\Source\lcd_driver.v(132)
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .SR_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .SR_SYNC = 1'b1;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/r_lcd_rgb[0]~FF_frt_4 .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0  (.D(n6308), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0_q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true", INIT_VALUE=1'b0 */ ;   // C:/Users/Yuanbing Ouyang/Desktop/xidianFPGA/T35/scale/01efx_bilinear_scaler_hdmi/ar0135_dvp_lvds/Efinity\ip/afifo_buf\afifo_buf.v(133)
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .CLK_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .CE_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .SR_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .D_POLARITY = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .SR_SYNC = 1'b1;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .SR_VALUE = 1'b0;
    defparam \u_afifo_buf/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF_frt_0 .SR_SYNC_PRIORITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_36cae626_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_36cae626_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_36cae626_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_36cae626_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_36cae626_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_36cae626_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_1_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_16_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_16_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_16_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_16_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_16_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_16_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_16_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__16_1_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__1_16_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__16_1_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__16_1_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__16_1_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__16_1_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__16_1_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__16_1_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_36cae626__16_1_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_MULT_36cae626_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_MULT_36cae626_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_MULT_36cae626_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_MULT_36cae626_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_36cae626_207
// module not written out since it is a black box. 
//

